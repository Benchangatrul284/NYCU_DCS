`define CYCLE_TIME 5.0

module PATTERN(
    // Input signals
	clk,
	rst_n,
    in_valid,
	target_product,
    // Output signals
    out_valid,
	ten,
	five,
	one,
	run_out_ing,
	// AHB-interconnect input signals
	ready_refri,
	ready_kitch,
	// AHB-interconnect output signals
	valid_refri,
	valid_kitch,
	product_out,
	number_out
);
//================================================================
// wire & registers 
//================================================================

output logic clk, rst_n ;
output logic in_valid ;
output logic [11:0] target_product ;
output logic ready_refri ;
output logic ready_kitch ;
input logic out_valid ;
input logic [3:0] ten ;
input logic five ;
input logic [2:0] one ;
input logic run_out_ing ;
input logic valid_refri ;
input logic valid_kitch ;
input logic product_out ;
input logic [5:0] number_out ; 


logic [11:0] pat_target_product ;
logic [6:0]  pat_peach      ;
logic [6:0]  pat_apple      ;
logic [6:0]  pat_fried_rice ;
logic [6:0]  pat_nugget     ;
logic [2:0]  peach_num      ;
logic [2:0]  apple_num      ;
logic [2:0]  fried_rice_num ;
logic [2:0]  nugget_num     ;
logic [3:0]  golden_ten     ;
logic        golden_five    ;
logic [2:0]  golden_one     ;
logic        golden_no_ing  ;
logic [19:0] golden_refri [0:1] ;
logic [19:0] golden_kitch [0:1] ;
logic peach_not_en, apple_not_en, rice_not_en, nugget_not_en ;
logic [6:0]  total_price ;
//================================================================
// parameters & integer
//================================================================
integer PATNUM = 100000 ;
integer SEED   = 5483 ;
integer input_file,output_file;
integer i, j, k;

integer check_count ;
integer patcount;
integer pat_pointer ;
integer pat_delay;
integer lat, latency;
integer CYCLE = `CYCLE_TIME;

always	#(CYCLE/2.0) clk = ~clk;
initial	clk = 0;


//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
e+Y7YO4XuTWmXKz1GjJTnb7ZAMKburbCzAE+Wa8X+PYEiEC6R5bf1Er/WzXNEluo
ynimjY61ikLauyuFIxg8u7S0Bo5EjWOr1yH2OX8Ab/fMKCI/1krO802eq+9KtX9j
Ruuca9UjjfByiBUCys1nPcNqGmAAD68PKFKsyOajdyBnVut6+95ZzC27sck9wIXd
BLX+/gCxjIh676jbr8xB+He9+nbNKpUEAfPZQToKL4qLO8BGqJl+StnPhYi8GtRO
BCqLCScLfY8xhhh8jnHTBsWEBqiXFNBcxOZp2dpCiYKP0UlctKK/wQotRVCfpYfy
r1wu01RjWY3ybNAVsc/JSg==
//pragma protect end_key_block
//pragma protect digest_block
LrpZfyXEDmu0v3O5YKyiIsJ9nMQ=
//pragma protect end_digest_block
//pragma protect data_block
OIHthPFNTcX1IOxsGlVw1oe4Ayh9dUmkhXuO4WlhjG8C9D0q1HG6V3zwDFkPnPbH
p8gDlB0PWiQcU4I2Xco5dU1hhFLYr87ovmBNa8ukvq7OyIR10k/ZUoqcllBdo1in
ezIlDEkhTvs7UKWSDPKgLUns+xH8H1cujL+7HQawPDJOTE0T/HwKd/TdlIlmFNXW
Wcl/jDYeYbXWRLtAFLGlBcvYpU8joUYTSZlkhFZ1/B5h2sULrSY+BIIKxrFYI5sh
V4AlY5qCUHd3dqJMUWsudGHK84nLq0ntre8ODYlR5ttf0/7HBpEbUh6uhoWd90s2
c6uWcF64I+59ah1ClbA7sWCx7k2PopkChYIAmuwpzqywRooi2lv3pStIO1XkoAOv
aC9uwrPux1+RqzYwwHKO5U2eL+fQHqeR0NVAd5zAfjYHrafxYAwuM24zAlguxD9f
gbQJqKVIdM03JWdqwSzmE2pRAXGnKX/U/E3uf3MeiVtbk0Hg9AGXdXEXzAWFvUXf
OzDjwEw32lVhitvTQn6LJSw+z2EjUFDB9fXWCejwu0Zb81h0cUFnyvw+7ZWugH13
aKRVPPkNWKLz1X2IZxp4sYtPfq6YSezUZ8Vw1ZBbHcFKwUjqoCRvwz2tDz0XvMyg
7aL9qI1nrCLYE18krdQbpufqj0e3oJKwAFL+ntASwf73dugBzn/f55mBwmFl+9Fp
sgX3qpZ50xVyRKzbfuNj3Q41Zr7yug7mFPa6lXi0Ahw7Hr14Zn44DEl3RBQEcZep
jF7GCihHMzGXBG0+IARE+gEGbOrDjgKIHmKAM9lh/yNClHg7DxS3Y1eHKth2mbsp
2w+5V5btBFSrTml+U5w0+Bvy2JX3xD/KWZnENjkpWTRdqGYE+IBBR3fvZK7T0rRe
Y+4GgxAmXBoMpj48vZNfzi7owMKISwNGbIgKNCJtF4RDhEr3tpyCerSvI9AN3v3H
NkjZnZdNTGYcI/ETMdIa3ZXPzSAnpdWDUyhhz4Qj6Q/lzp/eTzif8x2qNYOSwvrg
WYZMe+0zVRhvmGdJU9WFnVv2ohsk5qWqRJqxw6boW4EJZuWaQpUxDo8F2rjLMV9y
6wwomxoaxpd7dapEK/S0bv/AOW3/bJuWWH/PcLPCCkwh3BOwhufGVOkbJH4CQfBm
TaKBaMKI8ZbhH0/kxba1aO2tdmZKHv8iCyqkNjRFTaIIIvbezeuLmD6cfThleHyk
gVICIYMissssWHrWeGIYlr8Fl6xO6i4bN5hnIwoZjSqpESkN9SaGgQO7LHLP8+3o
cTDGJxNE43lgWqfRyVJNgexyrPr3RVIalhw2aN1XNGBKaiG6j0tyCORw4GhdPDmr
pQFQTS5AescR3l6HNGvQIsJSOhBBr/nU16/sRljh4wwHc1xYdMy5E7/f28FObVPg
vhTGG0mwiU6WnD7yyiNWBfHhZ3/50D3vWUHpfcDXLmwSFlXzxke+ecVyGr1a8DU0
NewieFcxbpgpHd6i98vsWV1RccFhddABAsdYlgMzIN/jZb1Q3WRm+ijZ0gpoJePw
rSx1u1ss2bY3LA6rElvxgJfmbKCWX5AuPPBNC9/xh20Jr4AI59Z3EyV76Y+z+Bd0
12Dq/2TOY92DSEEAVefEP9KmW4Zj1eQOUquQp3stbPwiVZMlS8SLMcmwChAnhT5D
WoxqO45uRLbQ/xf2wWmD5WqlhiayRTLM8EGJqUNWAJl6zHZhtBCpKq7zw5lHvl3q
tIslb/Wt+FNkunhuUfTxnPsOlo+umdBQoW/xKAlhmQlTb91gIvRLrdZJuu7uhD0Q
oDzwouPz/Rhb622YHRCVSueHcpnsDtA0hoOz7RaM7ZrQhDTTkrWF2UjOgRRJ3vRJ
hMqmbK9cvc+ae5P19YfmiciZ80wKTSPmiQlvFA4PfO6782ZsSUW9FGcn8BLj1AR2
TCW8cn18m53mtgfjiwZkqtb6CxH/41HhpSivpjk/nkk8jmh2P7gFaTRTvq+IMbBl
DQT+KOfd7JYfAkjKXv9SX+Ge+ICPgHnW8Py3XaRcAnCyNA+I/DmhQOT3B642Axum
1uoeTOzvgwettd8e+EF3II9kphQXoEp9iaMj10FUqvmRqFaNXBPSeZUJ8SyYQ3+h
G9RhrHU8IjRuxadaQ7AUTTL1sZYury0RG9BG1FG6QiArEAcHUsea5iEvEUpL8/3N
7+o08eVUdhMez6nj+ZBDxapEDLxf1VKAMOOaACZoc2iGZlS8u0B6Sl4Mw1/TnOo5
mpve7a0QfF+RBonTmO2INqhXZakz7YXGteqzjZzcB8aQw2ktzjGO3LMlYpd/kUgZ
JHVJnUy0g2AlB7u1etgnCOc9TAwJpFu3L8jRiKchmoYONERFOrsvMWQTjAFhuU4Q
Rc8y+X9aQXgcXjDHnSqx6xIsguw6p+PYa4/egr0yKeavg9VM8mhrdYN81Cpme6ET
DQUgp78ecB0joQUZXC2dNnYQoWtsOMLxSfRFjWK6r/2PTuQX4UQNtrmPotZuSwOy
TPejAJzLENbFCZW/lvfOTe7OKM/V0zRWJ6V/rYBJB71Tpc4XeAmr/A54zGBFxWqp
W8dbL3MNknMmXNRXfhtz1TGdEo1FzCEqfmaDzM7CHx5VG749TT/nRcsTObzmItnG
CW8vIMqKgNVxd0IyAwy03lfdmZRPhM87mJLa5xzja4v9c0Hq7HuHOetPPqN6Q2Ff
yDRNEN8U7klPoYP3pIcnOGoEHLonqlKCYw9XL8nVTFNUbb/qox+/knbJmHTnWuf/
tR0RlCTXRBuv6uezixH/fzG4UfgOGcPeHvfuToUPtOrBMOAbpoczqeyYyI2JiHgD
2Q8kXanUcy8KLrd5xgB0iKg0uh9JmFCciJBd1PQpD6dR9RCiXzxlrCA+ZXjxpNio
HtJ2I5L1WPbbJZY0AXjFFQKOKbT+OAUi5eFBU78JXTAm5NJpH32iiXCwB1P/IZU9
EHDF9ltX60aITdYSZuP7Qrx0MDXhY/OfyclYv1szdj2Ik7Lt3y2ov6SyYCcZODS0
81upvxvmYFOT/rccULuf8ZSh8UzNrqUlImo2wPXNpd2/fwwZCpHHsTDEeIC8cdtm
zP5rdwtTgI3cAEliOb4A2eqBCM7ExkyP6OGnHz7ul8Gk5QqlHSXloz9afarfKN8x
AzWfH7+azQmGttV/b5okeuiL+ADuuzibmtnfc2vfKsZe1VgEMdftMMpMj6pHtkX6
aP5sNcNblHMayRXe73ULcLsmoSR7W4LZtEEtomaKFJEbX0kmbjjV0YhkhgsAPNqd
fUnDxegXmSq6J3dNTz7YCCCXb863yz8j6+tG1n0rZ8RTIp5sgTkDHyXN8ZFvQpEc
/HvlpMQzr/AAhK2kIAE4cd6V3P4TKYzHnR858+cCQyOz8KCsCAeXI1yuLUSv8DHj
AmdKQ4rEQiczQkbPah0qz6S3Xlf16ooqrn3Tbmo9+FDdYvwadPNYSG7hcuLvH62B
Rjogg2NbVZS1hZ83MhBkSdeYDP1FXKzKIpwAaCVe30iFSfVUFOe8UiLQHYcVxNOT
3fSapQhcQZibMj97cqNctlIN5AFrf+B7+nH/q4tsSAlfz0RGTdzfXhrGrLP40nBj
E92XhtO6G0E98tvA37ZgNcAyUvSxvdAZtgxJaHpef8PbJlPdvHVM/s6/GMX2N8Be
vSBh3w/tpE22Uti651429mKau1XkErHlLN7R/QnbkymDZLNKdR6qTn64YWvEtHgC
iqKEmf1glRyUNbzQUCBDGClnX+OgTeLe4GQv+7yKQUyH5PYCGbm1kyEUgOsbOl/g
JmzxMr1gkEV6it/ffITN52tXD3eyls4lhlufTyPM/aMZQK5ezl0g9LfiWnmK/9Rc
UPjLBOKP+WwyFcrxrRyjAw+j57cUKIsFQmx7vcKB7aR6jybnrH+dKPbje+9bmQwG
yS1lyI7HUKPBo7Wx0IIV5TX6OX52ILqQ+NMVuSBM8fLerNDX7xJAVFh4rTrBfE8l
KwgIEXFE8pyOh+wtGQ0YHv8tDglvdNrTSwvNwt0ua7NE5WLT1Wyh6YSbJpm2DPMD
IYoomRe2btdKj8bmNT7MOhDS9/pErFkS9GUmDCdsxwKPEE3rtzYhu6rhDvdvHBdU
hzwWSWrBrRXzb0HrDRdqu+CUQRSms4OEkqkkRCsmelCxdOXlcHE04eyxU4LYgRS3
KnUnxSSuVFLQP7nasMrtma6bEgWuu5d6O5FGL43ewwBoc91MlKTkQ2jBgI+YaMw3
1jGp7o3UZ/J93wBvnv0fk0N3TAR8ncl6VKZBcRwhZBIifpSU6FQM/+xok2Z++Z//
uR8R6S0SEvR7qgquTnEY2E9rWR2h0DxAPukdV3Y2LEjVieqzLmAr7fdCTdZfGue3
n4TqyRFSRtf2edZCRWUBWT8GIo5n1MnapI6zMeBjXT0KvNIcopsU8CiAPEhv/xBC
TtukzMb9Dnz/fYlVX36dw7ilqF36mYA6SbETAGOI/H9vtkCooi4IEyZi5mOYqeAw
9vgSxS2r0Bq4unSfbtMHgJW/dfMLSI/lc7UUFRINuinTMCdh68xzs52mvZ5P9lck
r4xyhCu17cn7B7ZBOun57TqND35xKONkKZ9lpVChlhKVFZyVaE24MbRSZua9N7NG
xPDCtY+MlQg9XBVocW0EdV+F6Fu70NgZDnJzcIzBKa7B7iaEawItTj6qnhs4+CIn
h6bI4X7jtbi20rJkfhSQcPPK9Ep88np3qeBvT41nVWZDb/S+8wIk4wRiEazsEdRo
WcUjvwp1mYZxPzn2o758WIqhZVsVAxsU/8CYaDFHmfNcgtiyfsDCP4p7/7m7UfVi
y0IEs0RS1YPtu0loeQ1OOTsHkn6xCMVou1da+3Ujtd6b2bsIqoKB1SeiSU4OAbub
U4PUNGkdJ4XZFRDl9fchCi1xEqSKG5dFhNR5mz/WNcq4/z9QvTgoE0rpYOTv4t9F
Irumo56pziREEzwBHi9M8NFWgB7rh0Wq0EJJXnNCpxSJlhSY6ihnD97MEEOwL730
nzyC/Oim1YB8eiqGlQyLk8jP7z7Sco+xruznklGLwQFzT89x8nGUm6vKG9mFc3VW
WJVk2SRhWT/h8NAjJyaSpFaV4uKLfkQingD8LGd0h3UuXbsz1y/Tu7HYrZjngKgO
k5hrUAnsvhWVNk9LZiNtMJrz5nOXGzjTWTq6t8lW50aAWfvTKmzl9aRQgKUfF6KL
hAYFtQtBIclogUim6ZhMi1KpnHHXjr5oB4vsRQqoPoAogGMrT243XX0vVxin9NWa
cnDaICDF6SzHr6mJJ4Krtz5nvhKpdlRJkBLqaJcPSUZYpAs+M6YGpyXpcnDUoAzv
g8Zyo1LA7pGCp2VB/Y1x6RUG5eH4cxK0Z+GTPBrwEX7oSf5R93EHSqeXiPI2lrta
to7MVxu+GSy8d+2nQIbI61j5xuXIaUYuwelmKg6kUuAvueT5iqup5COvJJJqudol
cGYqRCh2meoVpVYPRarO5nWZREu9FcrpdLxXjusYagjIpDlpAeIf2kpxuFshezzL
lAO5ClBefzTfZ4PpxtFlRQ8FVzD8dP/7lNRAm2HrWrCX5TcHoi2oVL0/8SbfwwG+
CMf4CsxBCrk/PXFr51sdu9kTyRacyalSAoHQx18FANIEIRpb6tC4jf8dXThbumVg
s+3Q0uqNiOTzkHBV3C/QrxoAhRby0QhYsHApY3DKo0qHx8l7cSHaQD2+tCHYXQ/4
6mzl43dN5/ZhHZSiBHHunmvdw8ZYhuOZdkqJaZN2sHqEiLQwr/Avx1NAtpAoc9Ra
3L9qCnm0t4SGxjhQetVDBrPAZ64uk8kAPU8lP7i0EFMm3DWjYAmF1mWmCWFr1Ny/
nf4pKbVIa4HkeZwyzawo/U/sGp5PVef7f1kJUk5OBK+KwNMvz05aNt92epg8LY8D
ni6gEPrIw+gyyyKZ7Jnzk8XXS4qrLYyFalxB1cxr1yoNoBu5tePlRQUfIKb5oari
ElDsDmUkHDTpuw0adBmFHbuonVP5tTsvT3Rwaxr5yE4U02GQ9RSLFptAp1MLmJPY
n/r9O3ZbXmkghMrHgu7wH4HnHSDBhBHqejN2Pa6JXQBHk16VZJwoZqWtq3989HPa
L2e313mwFH/gQw99XHff+ImZ7xt9WA4jYWVkQ9uO794YlHgsmMsfjcMZ4DdgyANz
YjjQSgN8L2AjTZK3yxCtzwgDb6ylR3riO40AWrjKm0gzNGyu3yn35EAz6/hoHqpC
9dgVFSoBwsD5Y/uahfrdd7kExIUJrZwkyObJ9ROYK0HdkJUgUj/kX5a1DB07Ih24
d7pMla8x2hakmILWWfGwvBnxB+RPBKG9RYUkXJgv3cr2xG6Uj1QyGawp+gO0wC90
PY7i96fFXCuc1hjkXKmgyBZvM74pQadlWTHnAXCeJ3+LUqcHzeHtZ2RWmoXHeeC8
3bNNEGwNykg5CZLTpExxSjrfn/KvfYstonDmgUrnGp/G4h3Ndi0yHPIWjkz4uUxo
o30DogZ8xBMPrnAKsvXiDVLxw0uLXCG7KW659m3XOMk/2rcWjYnHEi4DxmJxt70T
IzZxiirnmeTYFiOtgpH+AcUclM8CI7uIaZm/EGY4Q7Iz/2NWXnbphcvVYcX2kNwU
jfr4q9KeWrSIgn8PklAIpKtqZi9E8QCxslH4w+Jb0s/eV5L1A0JS2Fn3eg5rxRRs
ZGJ/f21z7GSfuITabd4qEJIda7braW626WNNgRmuA1mZW427IsypfgzrDFQdAzPY
zlrWxLD/kkNqZCzymfwBebBD2K+j+JGjf38+27d8h3X2x0p244LW0CrpdkkmukSe
IMTp/AoKtbR5x+TFy8lKz5O1GgjA2KgeK2Lv41fuFRm2MNt0uPQgaDCtyuoS3kvc
tmrlh7URxFkAoOSMUfdSnYUOTKvPmpPF0BFAT/xPuGntWLuNIZ5LPZceuA7cvNYo
q1RZ7UT0Bo9EUHN95xfZf8adQoumB1Zug44834aT3/klR06thtsqpfrnS20+yMDj
j5zX3C53sckSUj4BsCRcvPcBVwhEZkmfH1n6u5lZzWRWfeAGA4kdTDQ0eb00iWSr
FH3+rnugUORI7vvKkMP7CVOKlg2aYiK0Et1jRaBOcUf6gp1p7sWEwHzyAm5x5D9c
AJ3sW1tx3RZWpUh814QP/HoiJIT4SYaGoqS8oHYa5ONxjJBkGbxGe+LIj+F4EpXk
Vz95n1MjwNDg1ckfEu6JSD3TOPNC/8FN/c7tqCCTAGN6EN9ZwTjoMiL5et9c7grU
OXVthSLmoReaZv2X6ailGkY3qebRF8YK/jyrkZzyVtf+KhHTMkgDB2te+Kbux2+U
tlkvTYG5cME8yiTt5DmQzbBi5QDSEVDQo+ijQdfGJhkj+2sjWK6ZWhLId2mgjGLb
Y+22RNpjbudReFyAMvH/1+PA1UyY91xG01F3gmlXxE5UXBYPgEm47N/iU2NpyFzK
DixvOZA7UCKgxwOfMj5gzZBtDVqz1pYHR4FtngkFhgxNFUm9fbrnMib+HQZufg2M
yMpjapQUEzwbXYi8eAD9q6YObaLjLb65srUmymBOyV4eXJSM6ATgzbyijpzhFgJE
h7jdWnZL80LdQRbCanlvInEF0h66GCO4g63H848D6Hc7jQnRo5pZDqwXM70hbo/G
e80nqkhwW/2rhNqSOkt+4jXmW54Q5myklDgb+/o0qMZhL2Idiv6koHqRNecHJMM3
nWuSdF48pAPhz7RyzcB9zcBTcTKI2xGcJyJQlgTwSILALchLtrPhvUzbZEbehcpe
pOIgZLCOc7CL4ZTl7mzPEqWiT5AJvmORkFYt7YPtLMduskSNKQ9z7S9gD6ThzHGu
QaiT6pajocBTOsR0zromJ/WrmHAP0Jj8C+ajefuTc2K3icra/Ede97dlKLPYfdG+
re7eP5kueDGCc7KRCqddkechbpqYmLDFBlTe1kDet8EeUk2lvWeY04A4jhWGiemC
UXMlV6PUGbA5J6R4TGE4UFmE0XvdSu8joXNnXk5mG9rPZA7ooDdQoN/e82PhQmhk
zNwZijwwPe/pebmSHBI8A2KJUyC/DiFPmT96CJ/GWRO+1D+/DqQRjqyF3MUrw3hX
3OWdSWl9V9UBPId/+oaAH3KuSX92SwLQ5gwESkhTRtxEzSUKskWMjkMcn47X/rzx
VpzNY5nVKLilpq1MGfkAlUOyfBbnqJqZa7UJi4Dg9KH73mXjt+eiDaO+RjSxdOQL
8zHZteCbAJ6hWbUSPPAV2dNKiGUwGx3eeiP/UOYZSsBQNmg6vgya5HUUEskqbXVV
k0seHvKjEWGzuIDbYzfijhwF1foXWqc8jR/rpi2aSE+DC9p+KyserwzZZ6YKipib
V+VYEESdhW+SDpa/2deRcYRP3yUN96LaOIqL8wo9eXh+PTi3TZ/DMPkzvtEsjIWi
aicZOGHsZq4UbNr7ExRXQKm15wlW9cIY/EkHJi/pOCdvaopcQV7vcaFexloQsP6L
+gaEC2XvMfUJbvxk7cBx/7ziwel4ACjVCzzy4gVwF7rtSu4qEWngxoxT69+ndON0
Z3F/E5OxiznQ9J0knxaxWbqsVjb2sbCAHIfNtNyCi8NYgxsq4TtwcmXt2e/Z4pZO
vhRidEtNMewbheopDS5aIxpkDpgZQMwJN/eyfmaDKLuRrJE1+r3YwsMXWZ7/eKkI
XmE81/meqUc0S8t8IjWvPTcU9paKgYTdEa2VAax5JXBF1tKdfUc3/5IlHV7x3FEz
njdEaGKXaC/+F4KQmhCALU4j0IJTn8gAGqzKZoYVyiEBYEl+KOw4PEs9Dd8Tfeag
nmO1sas3gqA33+mpWjL8hCtNLJ4ufTal2s2pNsADH8lhlW+B7iKJgS5WZuWe8oDH
xMMWd+deAWgEWyhoILEo365W7DjhPvmhc5LqHD2X9o17WEAsw+NMAFQEXDzt7ONm
2SrJDESc24xIcwqr6GjM6MBN3QfOrs6zpEOQ3bj5ZqniAcqgL6Y1bE/8hFsMGemX
f9vvJwYjNIVKw0iXyras9GSYXqcDCf6dhZQrWrq8bz49gXidOqv5v89twnivbWQy
881yEUqaiaDzmolKoQDYIv/mre+B8M3ZCT+SAc9km6ujlJUJCa0aAusunPJrzn59
zSYRnZNnJHbhv2eyLk65ufHBOTwFUuoVMZcTrjr3uSzN/0gqI8gwnEnJQ9lPGKLK
3jCX/oiGxWUtGT+tBglTiMZd1WxdOfl7QFQDv2hvmyYmrwkXqqB6xhRauJ5vx3jx
7tXWsIZd5U+g8jC1g0gVSfn71vI41lMpEQ7Z9a3DX+XKVWDR7o1YMR2PSwU8em+9
y2qrfoM/8i1H665yyXzyYZUGydh9fdWP50S2o6gxrYZPJ5bSf+hvGs/qngPI8mHy
GLfslQB297KM1e46w4KH7aXX5NcgpmdCFGa2C7b4LNuiIHrI6YwDAQS4c43Grhb5
WIou0+zZAt9Z4HMvg6rSbgaoTC10JQIinPWIlKyITyEZ/Eu4XtJy5y2X9/ZiLBJG
UiDvAy65HK+Gkb8ATXxGOjP0Ffv3ChDO7g3TDcYf+kaxipOPlPksyzfJb3Ukzlpd
SCIgw9ZV+eqkyoamOR3IuydjzZWUaVCdAO9CyMQZgHm1sBjyLszSlVU91eBg9Pir
7UMvO9NP1NCOb9W31dfKMFS7Qv1C+pkiOVGyTQkh+oD5K31Ei5fUY3Ca2P01LEPo
60hUaZrfyjn92UIK/NWsialsEqY2Xf+2lSB2/ffrtnHuSFmmX/KJ60GcLkeNemy+
2hVuXGHp8ghttTy5eARd00dgc+i5VfBs1B3TQyMVubt0GncxV6KuzoLzqi/vxz8j
7xJsIN0p6yUeRkW6Z962Qs/QVRMGWN3crR+eQu28MihZt1ew8tAakT3TXMC+D5nR
6HOCFF+lLI+cEC3s/CJw7dLT6ZSQ21Wnwagc+oqNxzjvricDsN6A9hxZRP8ESNEp
Y0jVaxG1/msKnnKqg9y0q3uOWdwfZO1z1PM1wf6kwLrFlu3oSMuHQo2C7A1trb+h
HwSar7nMrfeCH9dvykNwMeL7U9wW57XhEFR7YGfqKLENxJB6Xun1Q+6o2g/c3sC1
8/8FVo0/nHTYh9a7KD3aU71H9MIM86JIZBj58u/ieQWMHcavgJcroeRtBGLfJaAJ
mGsgOBwgL1qe5nyFZJb27NGf0rvTjAOEhfcY3bzDAQ9f9q4vonL6tprkB1v3Vbv/
7gf0lPZnICsKu4UVUkBMlPw8lGctR9jvsWqEPiXVH82BN6qiiWoBcdpQTWF1itMs
nDwpiSU4hud8YhI5XzY7IY+RhshK3K/gzRpFrRRQD5tZxo3OpFe8A5B0tjuxiHXN
nefAGxUHOgEG3S+OwBpyCHKvKKVo4oXtI8Q++SpI3d6LrxjW8u47/sZXEXt6ebs4
p3s9e599iH8/vwt+qopjJMzEHO2vbaiAmT+Y+UqHAoa+PZtntkjAv0ITRAkxou+2
7ZW8MIOY2nWhzT8EZxcs6qXF1KWkPymgSaZnMVF+6ptNGJ7FV5DGZBIQQNbd9sfZ
vSPanzI2AoqhXgxm1YAJ47HbGSPMZa5eQfE7TWy/3eyHg0nhxYEMjVquB8OBPuFA
UDOlYX8Wwx8Hs4CqMK2KZ5HKJWGfBZOIPW4rvayOP3QOqaWrhr51aU0nvwjLZeCm
kcwufYU60lj7hcPNTrB1S2qQbt07+F20V77pkhrzAwBXiF7qQ5fDyVn7DVnFQc/z
HKLQGoj+/xm908Nd8NFyoX3Ii+r3Sk/MlOFJbN8FbArm6yVJPf3/pDUunNvZGeUu
yxkzHnEBBbN6h6x3zVNCEPkxsach/NKiLsHKs6TjFrm/mUoNuj6+QZXTdniyLUqy
EfU/s2adR9OmEso346zFSLcyh4bBNd3xM69XV8OwKFfeCsqNnEVb3tA8LvxrbNpo
jQveS5GFNSnBDdGpv49ucIeVpw+uuGlNCrCole4dcNpYyEIeF+lDzo8PY5IQ1yh8
taNJ/TtL0EjJrgOey5gRufAXE04LKRqab2IpayYf8N1L58VZN5k/J4IC6ynuFyiS
q/BeXmoiq9bcIwbotaH2Y5QYCssD5pdQyKMm6YPaCdkg4V4bOI6GgL5yqYKBxzNb
8gljNTQUEP9NhlFvv8MtI7F9cJsHR9eVR/+qzagqf3qgCBI0fq8j/1w0BOqSCEy6
WeuL1uDr8VFytoE9HNUDb1QEOMhC7Xk0CxdEMtqnI/MS4kGF7mQtyH+wR7sEssdB
olCF7UjHZ8dC5ZADGgjzatBQ541mABffLG0G3OQPCwCBTlzGZpKLlgE69HfAZ2Q4
eBoaJTqnuua1+LmsPdyRCIL0uJjedXMV2FITdh3XpjiXQlUgsLuNpJxeuzNp5WRZ
r0AG7CeH8M2sbSwbDA1h4sWX0euk00cEu22R3a6TgxHZmcvTJmXeKzEhsI+Q+bTm
D9vV3l8ckKYd0iSsW2kb0jHvWNOurs1GWR7bnPhqRMviMQGIH6EYBiaIGrXCYche
e/BR3rgF59KdyqwNIODbbXgvyqkj947u1YRfOB7Z0bhP1q+RS/+Y4O+G3ZgIgfuA
VIOQ0xXkRbJJsL0AqkViL6L106NOWegBxMzAEGQuKclqw5i9JkKQifRSFNLlMGxN
OsLLtZW57bj7YnvFmHfsba+OK7UsH12QCUH9enM1EH5YkWyJHAGTO/o1c+u2VxCN
remxDeMDq64XR/SyPZcUEtwsfmuwNc8ibpJqejKLz52fiLepRVK2eckAuwE2O3Y+
d5wTsFijU62ye/B+DFfa0Q5lz91xJS1z6teCZOqM4bZMGdCTqHfUk3V0Bt/MHKAC
3Bn3A6FcQDa+MPg7XY0L/lsWRMGlLYUNg8B4GhxB9MNDaUPzDSkSq15AhZmhY2U9
droN883IsGE2He9LTIjkxbXzVaUwgNqEnGce7q4+01l/juV+jpTvnPbChiTAy+Kx
xxXHfSq+Sja7AQZxzUTOK7GEs86e9fWf2ebaNXQ2yN04qBJZ8NqkD+RYkJX624Xi
7Qahxw/u2oubv7oe0YU9hbgkjWlOyJAIITr0m7XO735+xXy/N6hu1GqvZ0l6K6Dg
m0idYiOv5T1MgDcsmiePBhSNAqdvIff2IflmTrZSYHRY1kYIPolnZO17bMf+ZlSS
JO9oYAo5mp10ky1bA33KspZfU0ozKQabwwXT6jHOTBeOGC0aO7KeDE8gco5tRF7w
dL1pHlJWx4UDwojNR+0gFdfC/bhtE6wir9RqwWVWMlEFfuo4v7PUQPADT/Ld3TRp
DMeBF/pZScf5lR4LAl+XoZViYa5UgIyJAK5qcDseN+IS6c0eS2h5hUqyPNNO+fLJ
0L9/DMqtbpqGyMS3BFQlmnkhRwvRysGeN/5nAIGJZdwRHkl2mDFw3KmBZoiNnmeW
HhgW6T39AEy4V2m8hozd0ttxnCAT8ZN81KnuScJnJcGw2eNA6Vs09js1ofMpwdEE
lc41uHTgvyLoGRiJU0eIwPOCtsuzjJWH1psULVYKSU5+Tw8/i+e7N5L0mYWs9Js3
Shqfc6oFBlKizFwOBjmkHBgI+QzHExjIPCRzwmV9qQDrN7cKm5n/EMchGoLaKSjs
ZEh1cLw/iwuJkwCJxgxeW+4lfkUa9x9XHxfIsDvo+sr0PW09vvhY7KQDXx+EvsLr
h9AbLyDo83dsOmWj4j4lxbSgW9FHrjjrfE+rJl3LLcN4255k/70ZYYibAVSfcItA
iacxtbm5rG9B7vGiTJLLvN2AnGoVC3t0uQU1j9/Or79VjiMwLTYXjxDOOEfuRRgI
jcJfYBqfqKGrsVcVr4I4q6EZg0HWYpMt2vn5Ci7eLHMNm54F2tEEYju9Sn6DNUyr
E9HXwIby6L6qGgRYUsUe6zwszTu0ZAsyEafxYs+WBf3v66trhbs5qFHsfiOsr0Cd
vLe3DP1N73zlNj3kOj61j25cKkhUTWXikgSfceZuwGw4oT/FKxik0gr1O8/ldmr0
auEDp3i7PHotCu8FN5t5oedmn2mh+f2GEjueA8YS+XcVIU5S1bcj+ZjEXeCegZ1t
wg5LwU8wYB4gV+PV0Be153gMT8FkNUui2f8F9DPdVfKfNHnYx/XTzfgt9WIU5KgU
4+BnBwSDJ2XWCwqW16zO3394XzzZuLLyCw1kDDkZDoak/3UdkxXRwH6H3A5OB/xE
Y1KlV070qYG/BETo/ZE/d1//+R3N7Y1ZR9+qhooxBh0ypg2Cxvj2i/1frhhIl//T
8OjJtF5o3+nEB1QG4/jeOxFVIQ1fd1ED02mVbqU0mG3r4FL41R/urAYZy/K4SXm8
bMa9pFoph+72X4TwZU3jnq4InWVyGmpEt+lrbdmk7jS9cf4OQybCdVmdN7D7SYAV
jREN6abux5VGXFmvF/q/TS0xS4m2+PFZqRWNw61XeapadIO8m6dHDzV7eNWcIb8/
45eFlS1OOqbJzS5hcz4TNnipEUoQm5/nFfAl4O12fjxJZYKCQJi6mJf1IgRu3w6l
Yv3wrX5wh0ehwIhqPeJm9CMAcJuZPlt9kGwowIus6RiK90DdBODLx96J78y55bNn
d+sy89/AxstJTALGZkE5oRKRagwtwdoWLIkYjVeNEKKAhWeTy8BzNjgY/IB9ddKw
8yzFyo+2J6HD6HfRxgoHbXnDezYHbgIhdYyvNtcuTtJus4+Fb5p8qfgq7RedCWft
y9slXWfVvMZFnP7gCDO8xRaHhmdmS08DVNXo9PS7JQ7z9WnztO8HeEXU7M/bFnJW
dbd45Nn8Vj3kc7s5x0qfATsQbuM0TQwdjF9spuiN+4BX0Pmm/4rsz+YIQzscuriC
Qf5XdtwU74ntWe6NJXbpmDCdvQizBogDzBwPt2qDOCJ7TiaJugV/Wsy/8409aXSi
TinRfNC3p2aYOoD1cWP/aF03J5mjilYhED77V4RAF1PBfFHhCAi4k8cNl4TbHeoe
qTHdEnyKj8gHEsJBa7zVm7ntiBPztnjSH2cjOH7aBCpZmXaQQsdWIPdYRt4LjN8T
JafbozqjWIpblQhjBv1nISE8AgiSs5S1nCwA1xk5dVk5FbocEUo9TbZKJODT6u5J
hsc6tXg6dpxsTJWDdQkYDBEjESciv66MdQ/0ekG6MRuLXR9uRXVPyArvU60DInex
16gPwZ45O1vMCtZJjMzyv+lsK3p8OCx3LW6be+PDyfw7I0hPyGP27oL978VcnA01
Wi5b/rJN29w4SOQ0gHPKphnCSVzfbsVcSVAehCYjLtyQP7JOtOCfIyONx7JRKGRQ
IRhAoWTYDrlzS6TlgKqlEpqPFUHm/AWvKng9mJuqM6TuuiClZt5D7GIDE91xJk+o
R13AdZKXGKb1TgYoekwZRuPgf6eeIJnZ8F0O0QdNwMrD5WUZ53Ca7rQd9J9OlBwv
k1bE8BrcAk/KGlmqJAv62sZn8g9piagE2JyD3fDUpX+QgUKrzGPVWGvhF8QGDK9y
Kdp+h7rEVB1KV+2uiq/O+izr/PqdO+kZhzYrJfGY6MUCDzz8lAgM6go73QOk6t5+
VHlKjB5a5ert5MEAg7Fl5/3sem29klBJPi25qs9O/P5qio3L5AMprHCBZ3M/rAys
rgPtzwAfbUdmPtxE1wiIY/do3NBAD4ZSFWZ1q4YfX1Kns4iiXDdaJdQxCsnlVM5s
kIMjRgYlwKwTVJr/Hf+7KUgS1GY+u3C/eYHrY8L3jvoDTNEk7wA9mlNyCEjdUm+j
Evgbv9ncJiwI4dHxVu4YlaFzDttiXH2cNTrLNArodJZLnC5HGK0jb0RRMi0JK7Bc
O29NFF2i9K/d20uXhRut95xotdlEgFpfXI2BBRROIG0RtcGZD6dwkCqrTb51ZrtQ
UYuLTLabpw5vR9Vt0gPvtyBMLE00wb1ncdjuX05xBy3hNtEe24XMwpuAsKR+w+7u
aT8MAh9fncI0lR35MuKOlsEyQi+r+3Gzn3R/ncNw9rSMQAtSAxVGr0hrc+wdDISM
lYYOW1bkiqtziuwbOTt6LyW/FL8wgfh1giZRvjK8IuJHxjglrwjrJVfl4iNHciHR
tb7f8EevWIdwNT+6jNvGgJMRJHMbaudaX7cQBcEqdC42oOG5QZ5NXbycTPis+Qpb
BbFwxr0L/Cb2S7KoB2Ljy2wm9/IS+ve8nRiOs4TLOtLH6HRYzNPOzJa7LEf6Wwt2
QAkslhmuTJMPsbbXXvitx+AjjKOFvbkvVquyYqemfkDM6xqNmm+7IKTcTT4Ziv8M
wuvd/XHYBsx5v58BM7AH+XZH82LVFanA4WOW0U94S6kj63npxwASDdSTjruojYiH
CzfC/nWyWEhubTZna4eZ23ncDewT13gXaNa1bygdaILDJYOCV4MFHfm0NL0qvoqq
7cTCthniwNqdPWfvnbXaA093IDR4YT7L6AryP5fXbEi4zhMF7ritZeVaaUqemUZL
n099Qnd+LS/7KhBvvc08cU0x03L7sHMa/isQqQCvxHylhhphiAEdKmBEaNlBhahO
YjFSXu13lRv9lxBhJIzK+9lZc2huEEsihkZ5HhHcl1qcmNptXu7o7lKzsLifQnj0
CnBNJ2QYB+p0PdBgkq+fzcoEm96lCeWm1nM1/apFuqKiDNa/0M2IkZXZolSaItDa
6aCYy1H5jYVVHVmPT6uiODghEBiYEJqGTfQsUyBJT85fmUPmSaiSgq/eENXU1PCs
0i+JWXSRlXegWrWlBJqAGAhph+ltHgR07DRFXFAbMMTSR9U2qby1NntiPnNSGdMM
vNam3NeZSQJUE+h88WcwIAwelTuyp4Hdzj/LzfnTYqfYyN6eswS/Imc4toTwPVXw
m9HnmIlXQm0RURTi3D3iPfv/NBqhpt1mSvRB4xBRq5IsVV1gdT6lQC/9hQCP8qCB
Gj8v2wKt531XfMg4zJU8IEKBw0rlR7EMRbRfBcQqSO2k8eEg23fhoAADV+BCv62K
GPgwadWPm6yi+NItTS5SDn0brCmBpkpJnFlYuzyDl5tyh6GvUz4rQ4/eGJiDE6Bv
jEZO5uvcAWzg4EUx/wdaHOH5nJ/+XEXc6r3GbnsEC7oRNv1gYNR1i4K/K4DUjqAY
tEyrjnhQEbIZIRJD3B7O56ByDDaSHxE+inltkH8V0kATeqi9+nMUTknOK2k/ROZS
Y8YxGdziAv8m5uGglX1OZLBwuTjNypKvm2h35qM+O4XLAQi2UpkBIfqW7zJ7B3/c
FVhX6hyem1bozfGz2uO7OFX8/Mnsj2tDnEAG65UxYNjaSXHnPQLGlcZwkaA3C1bA
HTcRS9Cx6Bb1V4hZ6BEybDO0c7O++Ju748wMwY28ESJxbCnY/9RFa7Qimp/gxMpR
99ZCejFg1a0WbgsB2P+oAB4FwEMo85QBBKc21+doCH8VLcvvdjiGciiX/ROp9CTY
OV5Fwr2qJx9fF3EcEe7Z2zeWb+tg2WovHOtJsV+e9M1D8LCmDYEjTFXPJxiaXQeX
UPxaqWn7VXQv04aROwieV6lC0wqWqmuaK4yI9e8n89+pe2ZNWiEJd4nrYc+Ar2Dz
Hc1oIbipt4WuyukjSVPpFCCK3atQqNWFyUEtIQoYevM/dMWbKPtdP6ZfPfJCPBYq
JpCzrbxmWj6iZ4j+XYy92i5uEYm6Ib+6S5yTmVLbR2zwvHof2J4B3xuPj/ZkoP9L
P6ymitQlUkifQ/TxQpJcu+q61i1n9OzWxBkQ6TBDnuJYbhGd0+mq4JYh+Cuus/Ek
uE8CAG8Bp/B5HlyU9+SL2jS+2qDmUov84bAtCm5nekYaN8v/tqIgVMNdurXRqRem
jzs7r3zKSkXiqlxcWXve+k+9bbntWzGrjeMw5iyAzfz5K58tjQicU9AXVg5CPaAG
1arUAknP4dxIdx6P+IWeSMrG5eZ9uAPONyXWJ0d8mTnn8c6zVEHvXuw1r/KhBqaN
+RKdH9K3IyHD0WdrvKPzyMIbx5p8JK+W6MZdRdXkL6qI33eqElOJLzT/1z7BNh10
etCfHY38yzDD/QYNOupme3wjdVkBJk9VboXcFXAk/37cjtC4tDUOZO55h9N9+ne0
esMD91bvLgi8UxbPV8BeGKEyiRHxLgm7+cj6cjo9qpApWZpr0kHz0uoKxcA469q+
GbsV2qpqyAQQF9LQCmvE3ggfkHJ/ghdR0Jh8IQ4y2hRFHgJnbGlJis1FJ43n+E1C
kX/qpWDVZXgWBlD/Kxcbdp3XwDNE4ADgmA8beO8nYi+dZ4beZTevlMCIHOg3rI7l
vdXrbWW6aJqMzsmaPFbwWQ7kuB0OifKEU+WpM4DeaHIi4BBiAEyVrbCcQcMCHKot
FgMZ8YDNUc2SDXI0U0rDgZiPRN3ZlMLM1aKtBlP8p2dA8THd57RqKbp5IJwANt0l
Lgw8kbcft6Sh/DiK+Lk32tcIJiuEVjDKpPpJogPrrgeDrzMnDAvvyGEcxhhOlxv0
2BGUI8D927WxUWeWKC9plQvm4VGL8FU4N3ZkclwuC81zu/9pSXcMFCSS6X4WS3ZD
p66GlbXyPaXA5N3BALdAVxgZJcK1mJ/1mRmDjaAb/FIDdnDW8DCAswUbDP5dTI/v
Bmck7ZSMR9qyqcUysxqZ+vMf4wAquDu4bNJgUmZZHPZs2uyhqwvIeb9nyGMvLqmy
gGYIo1uYHo+bp5Za2Kz8DaNwASuneuuSqPfJ8t1CXlCRGDvmmrsfVh4DombYRw0g
4JGkRlHtEN1KSgzn9NPvhWwVt2ZJl6RmkQl4qCXhpZvtagkqVIR3kpIjbLVoSZN5
4A03lES33/FI83wyLxE0lq2S6yhoffnW2Tpeu+2XhbMp35hyy6ZiY9WBE08YXx3h
ttnAs5NkodfEQ6WVUXXjjz2H5Z4Q5rcq1gZaPvgLGWx7VYkxNXcFYknwYYJLB8Pl
o5SlCgpa2P55r6XDlGgQwDRAsw3Wq8CTnlADvJLyQpEnSYd+TYPVV2OhffdaifKl
CnWeFGLTj/bIuWuOGSb22BAFb9L+kRDMcf2JvrprW9uWFsqlBZWqMS5SHqwIjAZv
m5rnygKxm01jNHO806fcdE2uLC95BcUOGNl/ZG4N31UmElwkRmdzbAm+AM30CkeG
u0wabNWi9A7bSPdHK0qk41DmE3bv9/NZas1DtdJ4G+44sqT44ZQo4lFlSPNuyjTk
3Azq5wYA4Amne0xJDi1d7LWsV3b/e48pRz/38t92gfy3HM73j9UY9OSDIGlRwARB
pR7cLTa5FpKc4WmeRpwTz/qUkL3sdC0mH6wWK2aIadToHXkr1EaUk8d1XOOo3L57
UspxcvwKB+MgygyLWdkUp9GKD3vnNptFN4LTsdCYYU3TOUuR1Ih5gWc34takfC7y
/gwzxoHwKtk3rJOA4Jv0542BOvVKRSvYuxQ5vW1hvvBsEHO0PvRiBs0la93rXOF5
XScr44SW9n9ZWHeoPFCeMkW2yDBEHN7afgqWpAHXC8gG8VBx/ktmhhIw/lA0Nrgn
9UUTt8AMJkx4pBiJyxG6RboNo4SOkUVjLi1y5l8uVJq9SOoKpVoIgQUOl1qLqKVT
O/OrJ+BNQC6Nl92Jw/gGTnlTvKM0UQpzqM36k+t5m9oDkqw2Bi0XM1Fmy9/lNxrd
KzhiHEvfFX9bp7xTYTec6AntQhEjqP4JQzdKNHDwZRnYca3tnFQlgQ+bOQKXD2uu
nLXsKT/LZvMf8M+m6YMkgY6Lu4T64tUIeScJdRBhfrzB9doYfjzRdDl5hs5uz/cx
T65PYGRxDYWZ5ASqHG0yDzEBUXbjzcDqfhkBY+P/D/LvAgIe/aMmoNMFp1I0aewS
tJNg4gvZnLj6ChsqKRUAl473MMLVfqyBv9If88WOBjDnWu/LM3ODmif8nrzhyNHp
aV+z5h13dQqEbB+Cy4FFZbvl0I0SivQmNfIgbGqhpDLIxIhJPrAdrPP6SopMlBbw
yRzN5biAnXzBVu8kg7tauohjBRItigpW/jLyybkRrWc4hwOu+6WsqYEdiBr4peFa
DAUpXEaW/YUfPJIwvezVuuRQ/l+9jADwv0J4SuVK+B1gM1iK3WnRSAICs54oZiIc
wL6I/pZbGrps7whLqs610p+X2xliO7cce3U9aHJmCYjF4gavRFq79tEB4H4o1rzG
+o6Zc5a/wrRjWgOibX6syFojTzlOn4N7ypJqdZq10ruKYtKKI2CgDrjlwveHQARp
vAh0BrN9j1njc13ekHHY+VwaQNVCtd2TGqGsWPR1T0lDYP2ems+qoPM13/X4YSY6
oTBRHf+XFciAs3ITImIukP95Wgx9/mrnycQk12ap1wkgml54to7rCP22JhitP96N
5ilUj1+divUcqvh2QcCn5iLvDaYVO5D6hsMYSYPMwM7nzqvWAwrpjYNx+hJuzzuY
3Jiz1ZOmGw+xTbvFl4HwEr0zX0U/rCA0lliS28/MUbwClA3m6h0AYq2rd1cP5v+5
h1zwgxZVnDs6Et6K91Sp5kMuBM9+Nu/N9VCE+Wys5mpKo012mcSL7wr+MnQtDolK
Xpz6N0ynLcJ22Tr4UPlw1PgFVWZDmau0nalUGOeBIKX7i9XJJjl1E53RRSVhQU8h
VRvnwiAoKtY0LOUtzHqI0Esw38Y5xXGUNrOFFE1KBBsHc7DSGaR1r8Cyp8FOhvQu
0v+piTAK1dLyLIsdf5Ri1abEUEoUVpZNYYSHxNNIuPgv7q3XhWyLxDyIGOW+ZDoT
5Dde4bYQYSVThiVJiJnSjZGroxYCk5mYePf2PDi47xc9Wje8fDtYWegOOfD1qHY4
BVPwppyquQ6iq0tXq3/b2jAFomA1ppoV3HPGJFRl+yIBPS2R4YS9mk5MPoZ4fy2B
TNuj6y+1rF4JJWCRhytGZwmCka2J8iK3qUxZNkIPn9Wsqv51vba6A/3j34+1Jskh
dBr4i3j5/FtkKZ4NovwiXepUBJ6h3MvCxcxFmvR5LtXujavBFJHY61I+uZ22uArL
ODji5SXkR2es2A/a+wmDs0H9lMWwfAYLIoNdF0P02tunrIJocnTLIYkwTU3ZMCcX
GtWSco5dV/YJMCQ1zzqZzXGqRyXyYs4jxQ5nvIDHNpStAWIIw2R4dg40bVxJ3HM6
O53toSptLR8BsEIsqah904F8StwN6UtfKJ70e+R1Z1j5aL64ozSzOkMFsSWBVB5/
ZXtAGfUdx9GhOJSZwUnTINVEPmfpctu8tOKMtD2vI8nMYkMkwPKojz5Q+r/HsVja
8bykvlZnAIQy+Z326MnlVaozgTfZixmg1PLGu5/hb47sLfYqitvA0vSm8GQ/t2S/
ujHAmx6xznXtJ1ldNBUHSN5mvoSpricQsoVzydfKPeWhFmn/gEt7DQvspeBzYDvK
ojJd4SFhJlkNy3hZRUYpQwH78wJinDo/wr8U+P7RRHHrFqiTo1tzmGjVlUvOoitH
v66ZcGYuvPCl6CtwlxhXJQguZo751IX1yTrdBw6qzsGAle1E5f1Wxwn0u7vwPMKG
Ki1rF2FgjiypzA6D6eBdFU1X5SQ8z9W2fNB2MF+W0DWxguG6daUXzhWNGuPinNO1
C4OeyO39k5GK6zg1megNa2tbVl4L5uReGRYlF1mSTbIhMgxwfTgL1BVHT7Gv9akr
J4ddmXZCvDpLdePCu9IK/C/NxslAMpk9irtsysx7ko85pznS/Y904oPopZfYRffw
VzRjYnnh35E+k4/Iw/Fc0hdWgUIPBz/3HOl+iqI6OGmsh9jDVf2IYXlWjeuxZBb6
rx+aKyCUMdQpXyyLs9Lwvi/pZGkjb76YJcDDvBloP+UVRdqnSzqsJGU4MH0xUD/L
6NsIV6zi37ieNDW6L3B4ACi2QKiDRMxkR5e0S9xsDRbL9zEHxZxrbhXK42CYioB8
zupB8pcdZP7S31628uMU2kiy7e1vsL914wHB3B9t6oMX3sZ1suYJcZTlN7pLH2Fv
iTYv6eRvglbx+AdAJCt+6B6FJKw7SB5dADFsIMBcEi5GkzbtCH2pyv+hhMG1Sq/g
eDs93OIwBni2caybEGuaZ4fGiJRB/2V7v7s9rMYYk3kEoYyqT8Be86KRCB0C0ROD
Bgza4722JV+SXH/raQCAOgKdk88U0k0au09sqWWQ6KOw12Y7f6Prkyssu6ALkPzQ
oIk2OdXRR2i/6AhYjhpCPHG0PmdsKhoopOdLs72V1Wfbhv+wm8D0P/dQtb5rZI3S
8dhOy5SE7BtWcO+hHZWRw5uWNAMESAsuN/PrXxqwMzxzOGW3j7GBIjB2PaZnD4Jf
8N3bNIdcEDZsXFvLMRJzrj914vpx13OdS/c6J7fOx2eDO/ypWTIaut8SIvbfjVkP
PgXwmxoGiVMswzDMwFqUb3mPM0E/dZ7sOxiBXo5GFzZO0WM14TVuqt5FEismYB5I
+YE+BxPLbcIffwSQ0qYUk+HJr/SKrW5kmrd6RpQfCCBCwgaXE0yNI4RE5sFAQqEL
0YS8C3ysq221aSxa2QkIL682cKRCQR6vCYpZ4gzOJ3E9HIvo2mfAORPgKsX9a2kl
zGK4gPfRIj5i8Hkl6/nkP7gOj83ZYylykELl2fJ3UbKL2TpXtwOmY4S9jKK52eNq
kuYJtd7b6LzaCrAZGT0w4Myc3vfXWDgrxImekqby5xK/Ykoaw6M7VuXcGJIHZwwx
MgF7XypwyuDeFKpPRvpc+5qnMxVqqvHn2uvMQ9KR7WfdBNThay5TIN+6WMl8EF5Q
PzA4eLfsLMX6/EZm/2aZ3n7sxWCFQK1f3mLw2tG4kFS6WFEEjDbKe4BpFIW70chm
acDp/l7rBw0cXnwL70J3DYsxbPRRg58GhbSU5CH2XLdnVQ5zErJFdvW+BFjlT/ux
xj6giSUAq4JAg80FHeWU5TKafgh2XffybkXqYWnR9GiEUkcFzaaueTdk1E6GuNlh
TGSUPeagoybVgD84zhHkIfwQubn/qJn2PwIhWPRGZLcH5IS6eDmZtY/rdntTsixZ
UDgqL3xr86BaKV2NpYbc3ocx0O6F79OizLU/ljmnCtjmAgywv7NhG9l6PFYIcPxE
3EgdH8KE1F1qxGkNrPrqDJ8aoKWvupCEl8b9ihtOltNDvvz5CAjCmzi2KsBuxCgn
1Wwg2YxL07OaAMKsOji0Ac1mDR46Uv+m0OuNHB6/LB+sSP5l1fD1q50amXk9pTEJ
aq//WmpXs6gGFuzeTLJBA23nFfdNCvsIxnUDgXToo5mu/c9JXDaidaJ9kBxCVY0k
1n52/hApNZ6OcUQgP5b6GwRAah/W3DYTpPZpNUdOm/lJHjeK+1U4qdQAlvbFXh67
Y/fmaseIKLedJswr1zrCc27uXaBTxyXP29TIEaXk97bT/4oC38r2SB4Ji42E5llO
3+1zYWtqs5GxvRqVWtBJt0ksyf/xH7ytG+xDsbWNOxei/2YKfuUdaeB0tNJM02nk
vpukKLXiDCuIGSppCrXdv2dDh5/MwyD1aczRPnwOBXlimwXTHlE1mirK3jSLsI2e
oMS8GDPeFsBY8rX+Cs0yYWtEJK2hqHLAxIrCmiM8ZmSCGP5bvOv5Y2KTdtSaZRBc
mr8MBb8BK8AXprgMzS3OYbRDEvnkRIS9GzFwpqcZsVUXk0fcUv3SrNhX4mhtITc9
DpJcbJuiqnEcW7VsHh1Ss+8U/njCZbmvsWSXetNJgTjiNAkhQKLgrLi8SDvTLpWq
o/wbMOyMM/nTUl0pQYhwybIklbMFiYVNufNhpVvVgAX71nla+dsilRuuq2fgbl+a
poowubgQYRpws58bCWUvqESf8RD2wmXpR2qdxuqkDlnmK2g1OuFBmyU3DxvCSbLn
VceCc4WX2tYBG5WhZCLTM9M+A3Te2Q+Wu/qO3ltq8N/CBYE6h+iD39pI8Fz8aGpM
EQDussqsXkInbs5Wi44HnC7x0J6X3gB6IjYWBisjDKxwEzKRn1RE8V+XlfAAcNfN
9Ao8kIjl7zUo0HNqamqMpBEjXKqbwm+SKQsJU5c3oupknlBlyRSSzeqKEMEyCDbp
3gm6jRNtyUN1Lcf3sfeldzPbAW2r+gjXQDkuOgrrDAQ8qhT7buk7YJF1n2uds/Qj
jAm/pDFdmViPVqvNAgATAXjPb3Avp+Ig1mE5r6+PbqCjwdCkIuMYnLXBydUvo59p
kSfX7ghOCZSWPdVr0SYrZ7qjFJwoOiovWdrV5tBRVoW6HoTDLUlgWyexkVbF7mvd
IWDpOCpnwthbrX8psowYBksSt2dhy7qHRHSALwbDQ2WS2EzqyeDdCPd5u9309Wck
hUFVR8qZefkJrYCsArrxgFReLgTj78n25DodOMzaHVqcUIMDoWLUNGXjHpvCKbAZ
+U6nXZWuZCdQbGQUZsnBuRe4/CVtvsA8R1uGTl7ppN5JNeVThi8WPlSZ0M5bHXiO
AqRW/jK6/t6H+Zfev1j3hLynp16ezw4J6LiIR6ka3cWPkHTXzd248/MHnl3gLJzN
9BDTHP5sjDWvZMOOYkB9pcLbfwSWVkzZybQTZo+jHxUGtu77OodymhUs1v79SANR
cxeul2vdqZiRe8Nj9JTsvl/zwK7vKsklcKFAC/oXMpZMGlUCHHq+EslDBxv3MH+s
HC7v9xptSSmaUCo/56USD3p2VwNYkYV6VqIgAJ9xcaVCwJ458x9ZqF0xtEjdObpC
ysY5Eo0y7HMfH9DRfo20ylD0qoAsWqigkRXN25smzSAighEj/SBY1xa5pALwAweK
pksOehEF4CuiinqoxFzJbT1ZUo0AXcG6D9UEayJ5fZCgKiUshfO5MxtfxzaH/iiW
OoRyT33l5ijBcMc4Lo0CtNROj3dYUn3tUVO+B8m68BZpWw2XfLznv2aTLT5heMOU
l6O2uwsheES0wi31AkSia9s4IlbvNLDsN6bMFND4+xawCAgNEt21LoWtZ5SAJVRB
xZvmxNszKJg+96IoYKSzfew0CuSrh+F2Bl6bqo1FUHarQ6WP3Qq9KFZFYcFXpT34
j37bZV3e9fbM7jZw/jcrYdPOKpSK9uILnKm2LXKnTBXUnmwP8oxSk+EZHTb1qOYN
Ur4XpYSr7NoY/O07yRc2UW4cwXeVQmCcwiDFUNq3sD2MmEidyILn91MfaItr7GG8
YjEbFR79PgmzaAY4nXRx1bMhU3pLxLr9N0pyZLfrwHtxRKjmpVUxFW9dWGiVE0L3
QrA3vF+n6p0C05fonunjaJ8UlLXcAJv5vS/2aZZQcawKDXZN3cKrYj7f3KaJBr+h
+3tQymq+Yo5PcKEMCUGR1ftPkCJaiV1Z/GXJQnnlJwgjAXoi55c3U9qiNPkJCfn/
nCwESmaEa8KQZnhI8+Ok1TksYkvNv4Y8l8B63rJ0xbcZmiTFs2uj/RJblKi/cGAo
cn1Ey9vmitBq6Ogln184oyCfoZzm+HOszyj+b8bZgEAjORpm39xsA4xdMGU2d2Cq
+JEs84LcmL2AL3+5yglJFrl993cPmsYBSi9vaVFv67bUSDeuQaiPUkv/+kvOb+oB
HWe8UeOqYMC7qrMMDas6Pz4+QUmBJ6G5x83PVsJzvcmMnLYCeb87GBWINzHqIzmx
PAUUcsMj7KzgkGIIPQonH7JIGYqVgzc7NK8Xe7AYSKySOHzBi/nzpW9IkeVVe4k0
4ELPHmsPB57Zg9LbeNcm5CWvxItmncnQdx0hHui19HgMJWbJUmu6BFAwV+9Bg3sw
/X9gse7TTuct7cA8znt56NDndOoa/vJo+sh/ge6Cn+LTpKgR3sGI5HF35iOB0u7b
Fe5udXMMQss3RcQHnV6sQgqalpmb2j1EVdGIeWd7ZFuwfvyP13Bh8zbJYF1zdl4I
yt//PZ1sMKN/7VRLdwzBPrXuFwV0nUgE4LegbosR/Zq/8xIN64Dedeyr28ZyY97v
OBgG/i2p2fqNzr7u7r7qMjztlqvA37zBUVhxy8O6ccCjtoiEEvFinBae12/DCQPa
dmGFeWHfN/jbI/5lvlzqhY4Nji64JP6HADo8cnGE08q7o5GuZehF+WbESMMB8YV7
oI4bRTpGfcQjhwXmSfHCLFuB+oB+kWcJRvCw0SVMLNKRRm+jONb0VJ0AQa7VF4fM
XovCyclzwMVnwkxf31jh6iSRdq6mZc7FptpOy1FbRIAm9/BGSyxu8Ykjo5UwfORu
BvyMMG5PAsir3l9Y+z8pXCApD2GX+BuqTU58BcMhjs2pDtMSd7vi9SlZ+acWTRsr
0EQHPcIHUlYJQT8cl0wXsQQD1gdj6N3LfIgoZtiSZY9vRz7hYI3LyAfUPXOMgsbO
vtjgsL4zlfiqyZxJXWZbOGxnQd3FR373fyPGO9/3jr9gL5cfS2cwXB9c6xR2W/g2
LVneYfXYo9XBqpnRTeJjxiBIzfPMB9N84C9nb2AVV4yVAC2gtY3rtzRS63OfhjnL
kkGeB261VIJuYIkkpVSZ1mcLftkQHfZmwRUmZZjWLGG6OgWowwkBwDr4SHXqbmxv
s7jy4XBARlSiUZ3fb9RV5wBZMGOixUNealFLm+rxD3eF4BT1CxBIEyi8Fm+Uwj9U
cLyJ2tllW5kZKoqKzuMQ1+ReQ54r8bI/fgLfE18qckEyh2v7F5Yzr3i0QNO80E0G
ccN4eM5zscT5MoVs9kIxebBEb59uj7o9a+AXRtVoDhNZU21TDi6sNKpryeSABH8Y
ikLrdhifgn6H9Hi7B8tcJIf1laSLYk2iWBtQPVM377V6zbbpW/ciRcj5Hb8Xlspy
LKP2KOQ5ojaB2D6N4yjsIAsfpnFsBw90gD9XuDnMMSuUYzrcoLOAvvsiZiJu5mrX
O/Q+EMi9Ebwm6jArOy4IJy1O7+g/h+5LDbQGiZwi2XZ8IDbpsCqfgkIlUsrAcVIS
ZfJDMK88I35+2Yun7AjgUQ1v8VzZe4legPCUi498wum/8L+AlIiVYpk0TralbSjz
UW3FS10a0todJwRRu5IGHgYexCY1bpq/BoKJru7DZZs8Hs0nlCY42Lno3ql9dsuy
rc5iKtQMd7lziVhyrk7yoUgCtKgzofMjeJ6JQtM6VBRHERBXHIkhAp/LwVjEurno
okXUNS0wwuW04L61hOaVvfAIFWqXbih7sqBx14A49eJkKF3CrwYGFW9MMCPPVcDz
CdDwiD3Zz6XhaHNsK6qOGg9qbGgUdEfz3XLqw08d3Ab8gB/mj6Lg3OKzGsnjvkg6
UDFK7NdN2ocla6FLoguOs4M0y8/FWAADZaFv4BLTmObIAK84hE5KcakyVw1w20Xi
FvDO9O/kGLCW6NexFy2k0+tYifrNtQzip5X8eRhYaxZkPgePpWrZubmLZMqPRg+h
AlkAhmkplJM6dki4VSU2XhydG3ipiUg2nKrqg/SM9dfUsKWJ5tQ7xXelr7DCCL78
Tueaz2wR3riiBj9HfAs7nU4q2H4IMSGukHkZ3JI3lZSDUvSuHNVOeNS6DwWtulXA
8TSvGbxoGUTN1p+7yM3IxHjMm8vXPZqSw5jQ0lUt4S48XnzbhFqpLe6LebK0y0f9
iBg2llDw186yRVgvZ3Eny0AHJVClZfzzH9IJhVP8XGOJWzaOpWLJk681QuDy8mXM
fD//FPK14sLJV6weEitE5qOq+Nd3Fk/OE1RA/wOjXpna2FTm/ARAvwxlQId4N5vk
UsdEFGzCMk/d5gCaVTRI0yaFs+iRH2OjhRB4tAanAI1XOZ//1Di+V3pVk1KysAqt
07dlWOKPeoNZDQvP43P7OICaw9hEsDsOecGWSvTPOzsib+ui8FMwPXS3bvcwyXDA
4lL0V9y5VbOChThF/LJtTXs6STqY/hMkaVSJW+APU8U79norLOitR4it5/0OMXQ1
uuaH8dN326ZQ72NxLTDFHOjRF74X9NGGQEKBoeMHwMMe6nPKeWTJSBf4cnDEgs3l
VIKnJ6TkeatJaWfv+rNIwWyrik6sVwYlwOeiCXtV5EFGN72jOuTHLJDOmlsl1RF9
h5Fkydi6dvpmNk9eFYi6bN2edaoSowabqNBuJuypYFhix3mabwUHcP5wzYYbTS5S
fsDinsWQQPv4RWOtuEyVQK1+mczpKI4YCD0Ru/rUPzfO16RVFkIHqTUc9y7fDN2b
FKqfEhR2NAoFDuGvYC9bgxbDHxYvFsayC08n+hcSKZUPisvOZ+fw5acAaWXrI3M8
ORjg62lX1CriF20NCG07HoHPAnHVP9paygwhDtwAhqDi8/2daBfklwP7FWmhztpI
lwSemjbFZdYhQqieQ5PI6/0bPWlDsLrncGCGRbE+lG1R1kCUtdRmgWG+7r112wb1
foDXkdyYSAd7Fc11RPXZCGtr4C0ke7RykpXxoQiwpBWuJYVyVuDbWG7cWOWpkgUr
n2Eorp4qgx//GAEvu/ZKodn50e1sF7JDmDnEvtlfx8eXMG0bLiyutTJAqH5DTQht
WOfLjSxuZfnMicYdexW5EwkGNJgLLHBVqBFV72e8gN6wNcI8slZpvdJKrG/2lEU8
JptNELBfilSZvc/rACyaRAq0q/5H618WVsjhiswqETVRlAAmGvjs44PyXW4amwrf
MvvDkr3bB1q7EMBwm2lTuC7oJ+6OIlAIDZ9iC7lKu03PHIW83Jo/H2Kp7q3pJWXb
Phst1WXvvutCHDfjECiNlInf2wbZQtZNMLoRofrya9I009kbUP+uFK7SdNfoIqaa
8YDGlkOjj+iHf2Iblse+/dyBfzgwEtPhLDoGTl8WjEzcVHXWjTVZVwgSsOlj7mOF
yJ6rsqhzeHIalFaL3ru7Eybe1uUzznRvQMDAObSNdrNA1kTKyiHUTy8uI7F/Fzfn
P4uLV3lNsJCCGz4PLG/hmHG8zyxqAZHQwJEkjDZrP2JQeRqMC8Xucx0mvdJGZ4ID
oSxzbHBkZfFBtSZvrq9oeQN51IIqdnSp+qvZpHXeQsPTvkveycJlXnZ8RC5q2U7S
qk941owXQx1TRKsq82D6WCsSjEcw+0Vbs5m0S3aal2EXEz33gaPck9OxHbetvSBY
NrV1rx/bVkFzSWX20mpAm55OPyzSoWa1+H8914FYtJohoZd7qIIpUAFfIZMevV7e
IIpW++4qEE1dbibmS6s2K6M3fx/K1+/MU8s+aiqRAoFE1juXZTWMusX34MUokeCo
fQgjG93MG+nbqTBI5Spgakl0/+BCNWFyUR7FfHeDy7UWMGjuhtSMa38pqOKeqFFd
TozxHJiTXPeaxwYXjt2X//OxFlJw+AghcHocJqzylT+h35An8nIfrUoa42DC2leB
rg1xnxNxC8hlrjMmj1jyaalxkIJX/hy2q08Qom+CWCK/VLjQ+T0V5cy5bI+9hZaZ
nfICEM6/S1MRwQ/s6HKJnLGBzGjQDN0KejAR2ToOxUr0ioE8sO1l9roQNYYh2xuW
aBgUBcTC+l8002KUfeQGb2CHZCFklR83UtkzTMs0sDKdz/Z4kFTj9fNPPDyY3A96
HPC+RdgdDG8C3smTGogpC8rqZRTyr3sMDTmYqA34SYpcOhaHSnHNhokNtWhBVy8k
c6b6DUTvbrqHLPFE58nBie5TkR6m64mc1EH+fSMq1BczWxX0dd8SXYMn3CgnlWXI
d96fv/px2OXs9cDkRPxwvA7eeAlhdM9Wsf54TERLk0sGjckWuLaIzyJgKIZx3qaX
pOiL3Sxg3NXuWhHvUmMKE+3z0MIc1WhO3b04YMoGCyQkB6naCYLfJQ/JybVjIw/F
P5WgINuwy1VhVnigokOHFB9x5cPpN5ewxz49ujjLbJgf933LzyRLYrngEYo2rsvr
wUpLoeYIEygV+IBBwDsOyYCIBzCGDR9imOwxXhFyGcQoiGQthgPM9HgZWknvvuAf
Bc7XWeSCJl+qtGBHSkFQRnKDPA32vxGrHnlkmg+spI5LMZ3iXCLILj7P2oJhG63P
+dwa+tyiobwyYgr3oJtRZi7UpveQY9RX/2Kh7c1D9DGERenwUJv/MZpbNW6XlOt8
aqsaeqo/H5t7ggvw4ZTz2bnYUfLveVM9/6ze6yoD6M6E4VSHi2uDhVjMIq4KASVB
Qqo6/us6f9hKRM14WyyeDSJkxhrc8EP9kzRTmgJ4OQTu8mUyydmp0ZF/NAc/78Yc
lzyRF9BMLgsdF+r5S+odfA1rljUvzcSHV9ojUSn7kIHHw0z6tmYaNGzMKFga2hNz
6wGwTfvdTABGKYrkfcrC670x+oXfVxjUMTmjsgv6n6T573/yRXw7VN2CGx1WShin
olK7E8R5iiuLrdV5BY+NEWbODtsWD2B8CAuQvr+hJPYCanS6eVrn9qfksmUTDoYG
pN9SGsRjEA2LthRjYJrG7SIgHrBBbgd4AMerjZ2gUz0hNzZP7DSUx4gaRi/4Rwis
d2AXXCG9qUhE9nriJM8fkUN7THqwdLwtZM7/j3l6MXpOdLhS22+blAtAKgMplJ06
DxilQvsdFjjE/Y0/QHq0rO5AP1pMQF7VgWP510Dtc6mjKvzd2mzGgIMCcFXAYLpq
yMlxgYzHEf8/MfGap38UJLyr7payVcY08gylsuiCw3nbIc2dawj9a0RJJ22pwlsQ
jmZFijnXQygRvUqeIfGceXLYIVAWDXvNfIn7elZNXDYdi36hBd83grtrZst/SnDd
+BxPJ8fQ/+5xXNaZwlystd2Pe8B00V/lritg14TN7tJ0U7RG3RzlRfDXWhRLgvc7
NI2O/IUjMjG4J97MRLF8ahlSsnNCFnYmC4yHwr4fDUWCs0zGVvKyiPWHXJqAEm76
YoY56kRMO/oiIHNsdoB+3Slr+rrzqK0Zbt3a2Cu3iRFm/Sc48Sehasa4woZh7bge
N/zKnAbTuS9deO3jzEbDwnm0A2PyES5lICiyi72grL2XZgBMevh+fwykBJzd+VZ1
6W7lqh6K8Q4mXK6GvzHWKBN78FpfbzTYYaGhmP8lZbb8XJjTYZ3EBeIaT6f9DDCe
I4Tn+UwrEuhWcdFbVHb/jBB1xKiWWWdHuAVdeqcCNfrlGZ49zuuFFq0iunX3urQI
4Eck9uAo6iukrYYJl+59zdFaJpGjynFdIJxm5d8BrHUNAR6DetRjSjk+lnlRbWhB
v2jrYNzK6BruYdR1cw0dnqp/AnVf5yVRTY81yaRuGWEz4Z3L+RGn+DD+1wwc5XaK
3b5k9H4e7X7oj+fdCa/jap/xrMyEa/W7TYFy5hBCUSbOpGgVfbBZ8ZRFGMKpA0AY
uQX9w4bKlVALL74ys/DeTNgtzKV05xmorNNhZgoJho6FHgdn0hNVsKY2fg7F9wVu
SfTBOdsxeH5RkRVOUXk1P769pRiDA2UZ5K/65qI/1MqfE65uD+MbJPHi3PUngv6C
16NuzDgwE9G0qoYK8MiNZqTUeNBvuaWW1wRYyBaY7uaLQuRZ2SepysdUIjTU8THC
9q4BzV3Ryqrpqk1CyG5PvpA89qM/SnWIOirDQciz/Dg1pN73GQasNUc0tq1KmAma
z1O7bP7tQX9jThcqfdeu6+7vROCttpJ/yoCyLu7/p8Ghuh2f4MJF3rRq+qCpnMl4
z/1DCPhZJ3rU/QzzA1ZTOtBDuycMdv+JhR1ymiLX/hBmUvb/Y78+BpKJCr9YacNN
Hob7SoWillcOApVQfSHIhoDcx2m9so38mYUUc+9dn1EWrnVHTwm8EzTDnzhlypjE
3JVqPSQbqC6wP3TYq1BPbTw7++yrQDq3PKO2r1IsStlrxQyII8vV28t+AIEixKc0
SLfGDAmQZzWvWvci50nuaE6MtRz9jNnF1xjVZ1qxWULIaEgDIXn5gCxrBa751Kd5
BdAMH3RvtPqvo9EH8QT3HHufxeP3+xlVNzB9zlz6jFDxmX8GMplFg6K5YGY2zUwL
xbVotDXNenXvRA+nsdCMwg7+0PKOpHR8ZRTyxW/hOFbtypBZcoZrJXuahhLlki48
sqwEI8jp8Nb1d+7DgtHeBPnuU2m/rSP5mysCS7vpmlT0Cm7UaxILj8BqNFgmhz5n
/JQ0yBXErpisDQMd1xkz1C4nxS5IM92B+JC/yuMLyUViBp4FZwI50chgp58MXMHD
cPPBnzWbp6fjeW46W+oe44DFO4v0HL+pQX+5y9ctg5sBOI9fUD+Ptfqi0JL0wKnp
y3tPVSRZi2wA4ydzB/NCHTROXJxkV7Un45XgT6uG1fRRUmXtviVgctXeF6zQmCua
CO4KEEUXYoiGAo8NFFkBzjV2FOrftNGRIh1wpXRjtZSsbsKKQlWi1BdD1e90mnyM
3mFUfC3tuLR9SZ6pSXFCVRKf6VOl5HywLXs0Hst5F9etKpZeT6/wpOnlqLPJq3T4
kXE+UFjlynPDVh2SBhNUXwCnrNtWpiJugD3IWWOH+EkS2ty4ybuNKiB5iKz7EM8L
7pXPhb1YlSRE5Q7h7afx56hjrcNRGeWjZI018K+jX/e5/wi9LRUwOI10L4Gyr7jP
mKevnYqZvjfrv2RMuYXpklWEF1uiJyEzVPC+w71jIoA5QKEeEPDAAS+V9ptd+SfC
8oUrLNWDCr2z9byWR6CB6Cxxu7sKPft7FY9uSaAHl4yhAvkAcvOFivD4+4ufOXPf
vAv8+nuL3lD5IRi2sqUNoxMzzDk8ExmoZZwHP5CgL+e+jU9wu94+4KxLSXqDvUUf
ZQYQaCUaGt4eIkpfRNT/X+tOIn7evdR8QVJMLLbdGcjsZY2bpG5iNB5CWGU8I5Nv
KG61XD6LfHQuzQeQvaFD+FCidcwXktPDbsMAIkL2ukskHxANoex8GKHBYnVmP1/L
WSGOhl1JBwgjW4v7efGZxpPa9MJ8WQ2TgfbDp0aUOno2Lg3OfaisPlTM/QcsX3DP
6tiXOTqVLoWhq09Gf0jFgnV486VvNvpOxLpBB02sdBtZcuM6gVq5vYTfOHoPES6t
9oi1UCkwQV9M+XtSbS2sze+4WaNe37N3Q2Y9N0xujjaRX8pI2Y9EMkuL88sRa6A/
17Q73zxImjEreVYNvtaYNLQAyZR8Eg7iyaNzn2QDRburmNKafrGQxyhDSeoT88qE
f0nz/kEr0JEx9AwEYVRipmoiV3cCl2sLjZx82t9WRXr6k3rjPtpZqQg5cSyPjJfa
o/qqWLE+96gxXky83WqZJzc/z++TnJfwIT3IcIWNJjPWW9rqIYI3vbfVAKIle7xI
RLzCWfOMsxNU0XbafW6REZRxOpiRUc27oU9Ll2yw0Una+OX8dNCNlSorN3PRpXZt
4/6F9KbX6VMHQ6U0yDcd/S8wjcstMwy5lK1WikivIY9z6xdWyfp7gbMN9n1Ib01r
W8kjwmf036sK3TkkLNWWu0nFd6Xuwp6t0HTXl+lW/R+YfFO4qS4kEI3kpxoApgUq
46kZykLk/s8GwABPMqcZCDWjjBe22flGhRub7LbFzMAnBI3iNuHuv/DiueYNEAJt
8yMg26m/CaOkVDvbMjuYs4YQpLoVqtW3MQ7NfF0tM0+7A8hGpYChhAHuEjJdD3FF
DvZ35HKYD8n0bHj2VH+WeCUtBMEZzOcILXZo1rxV55zq6e230vg1ocaFrP7sipBk
y6UwwLdHLk2QwiHXLWtVdMWA5phzCWLmFnHntgSStCLPpK1s8mMzFOdRJU7RQWu3
+LjAe10eNHOh72zuzNlGk5CjLfDl1cEjf+F3il7FiLSxkBGE/qrxnjQZYlRN+VMS
hppcVkUou4c4ob3N8o2tNldNMPnz7sfGV1E/8QfnosULFhg2bKAB+b1CMgcHBRlu
LFbWKSRdigyYtkpmcAXpTLD1k/KAvIjQ2cLbxPyStCH/gPXYnvqcROCBgv6Ass1J
i1qMp9DQwGgTTmg6QAbAeXmAzpYGMKPaWVMdhUgwgB5gcUl6UYTBrOSnQumZvMZA
9St1z9Xo8YwoPVO5O+sa5KGkPxRALnMqEq67glvcMl1JRDbmfPtmT6c+UGXrN8Mc
2vlr6GIcyw9V7oCsXkA7L1iSzW1Sy8JaIgx4r/4+jkwJkYMOPYlaEmdSt9tyMC1b
TkuAkTUBoFcv/1knE4Ter89joquoSwnTDvhUpKk1NKJdUI6GEvLF7QNtY5NmrX0m
nahVU7X40dM+xfkGos2a1WcxhPoOWQ4UBxAlK2up0yB/AK+GMyWUGHyjVkx7GDlN
3dL8X4C9nn1zINl1a0UQ6y+szabtwJXqbo9M/XnC8xeaiWAzdxS2+RhxEHdjnHpZ
1HekNdOiZXcjuJu9ZxSbLJcFAirfsfK78ccEthWd234A/5Mp97PJl45Cp6K5b7Yh
kiHCf0irWwj+BvlCyh11XPW1HOdXTySP4xS5ULrnIiEi3vksNL/aC1jRG5MCYXJG
SUOSHMNZp7p8/i0bU4kodycSZyf6b5k80fRL1LpwE8eHgkV9KMGBsUQf16CFLuKL
+TngMMhqy+mZBjW/61/lm0hZy0kSbBexXGthh4WOu7eQK1bD3kEJi4yZpgBffkF0
nQvM9JwRTS7/NHrjy95MSJKaHehnSYty5JcLNZ8cl6lv6a63YWKQmYfqtVxJleN+
w0UMTOgVcSGEAG4NQw/P84rDbUzDvdabmukUevuxK6INjpEjyJ1e9nh9qTAhxuic
uf6aAhRoX9HeHDyK4y6+LHxhXYHTQYJpZ/prIaQuM5Jo9MbDZ+6Hv1hfsusi2rbH
7kJ1dpvqJDN1lAJoXGOAUMknBRv0CNsN80wVUVr30/RB3QqevEERUx2ZanqKgQlZ
dDugfF7IOaPQH9q9aMYB0S4IkzkLXBwrLcerbrmta/TS676Nu/QxUCRX/BLeMsqG
Y/BnkAgVnHhy999+j/02Eee0BUEu+3dS5EpOcAJ4aapjS182arhYGzywqMvP83Pe
ACmUrHmVCGwdz7IdoFQdUtdsP2Dv0rkFJWIX+Rqex2APqqFBM1ArZltpzUlavePZ
FFPqxYnrXnwkA0QKuvb4UEh2T9Z76JJ60KYwwOG4oUrlUotu4T3W5CdskfHjSsML
WY7AKI6+qWM8ZXwC9J3ecXA928nasz/AhtczbwKr8Lrtxt1gsOHLbPA6bikk6Vm0
yACNkwrbpnDn1Gxiozlc+B3OObwVCuNsJFc5UmQ104jmag6oY09iRU8Gp57uYRQt
jWwPSDQw/ISJSMyXGoWb5+OB7NtjGlfGhE6jMf66INzzzu8pBxoTWIFNDW+mqwPb
fdyeCTzHxLqCfL3swcs3HbyzAtu5MtUiDm/oxA21EdW3vs0RB54M9qOb8L7zlCBZ
PHOucwy97564K+WCxEj5NLQH9a7EdMrWj9iY9mJdBGpuhI4QysNh+MpJrSc24fJj
vDk1zMwJ+4rnbEYhIIINpCRO+6jCqrx3WvK40gB4GC9ZcfQNF/lkcYGWm/k+jtU8
I6p9Zef9e+YnbBhNgKU82Qmxtkq47H1ZQhFa4bgZrvUGBt6W/CDQ15g2XP3dXnVM
KsxjhU2SzoPT86ukX8bmtylMeC6xmtAeadzhuguzs7EAYbc17bTVcmx5d1yh/xKB
CQufjPB0wqaBx3JuttpTCjKzmhyluCEgsgg41vrQ5SiXZDn4abrcNE88afNaAASH
jxOqAST7PpnnEpbgal/0LlFYfEQc7gcdjR3vADGzeDjHab8+F4sdrsZgSzPw9ox4
By1NxMrjvGqOG73XPYke6gXt8PU0PwcS/K1J+Bio/2os3Kfz4ovR4T0+gLoVG5Ou
mP0BnfiHl3ZKsJTgS+nOvvxwLVERM+O7N0aUbjNBJzeRHFsYs6nE0E4l1tHDgoUg
u8Rhg7O827re+/rDlz953uGJ8RR6GlsYf580oyAV/KLn9z867fYUxwhIQZ2vVAUD
wc28/wiNzs2U4WMF9SJ7aWbwkh5GR71A8vMnlHbVX9lSDR/pm6Ii4AvYX12deiNv
BBOJfpqkrYM9p7sJJtTyLLS+GS/wpSB11/CsEYbR/S+QymJZByXN94TrzC22Nhex
yH/u0jwxJLwEzs3ng49/sQ+Wax+okD+jrx45dR6jOyW06FWGeSzVjqycprC4oB03
CzhH7P++kiBEGK5FLPrUNS8zEgsWMn+u7AuoCAs+dDCNGdwnOGmdPaBV+zrE0Zir
SN+1a4EbghqFYJbl8rTSKYFX/9Um4/XFGDJIjLMmk8oXQk6QTNN11Wnzpae0adBd
s2fq0XbxCeahVyr1WWp67svy7ppZJ6ZPkG8kxj1voaWuuuzRnudxucSbHNsJJ1pz
rr5Y2K/6hQNYg0O7G6Mo0XXEVmjfn3djsEcLqeojdn5H2DPKvXUT98qiXZJrm1cU
/+MZ8CY3WxS1MCtU9B3vT67K36JT2C5PFQXIsw2S265hcOceWza6FhYNogrbaFLT
a9jR6ao8oQpRscjQW+V8bhWQ6fXJIvryHQB5ipcyQgfSkV9mv36tdpuk8VPLd/j5
qq4NzHCcBRtnmLv36YMAXupWPMT3a+Zi+lh6rFVADQqG2vhAqgFtLj/Xa2MWH0+R
s7+1JTCeX9a+bDdRtoRa+vbivy/IDzijdzFFslLvxX/uVOIg3pLk3PcOP+jB7IJe
Z1VHoFBwWMeUW4N37pJbPIoNoqDRafsTWK0xDs6uVYJpTIu2F7SMmSjEu8JbXueW
Q3XqV8YjLsyKnUM8xzqTVPX2UulfIDPPZzvWnXywC7mMLaSc6uotTWZYMu+oim3E
TQzeqFX3ii7qTXYL++jQuMEz6II5duKUFRYdgaRiW8mofzrLPdGuX1kXg19HvElK
GI1NGFEkB5nd1Bf/t1SJMFo0PxgbpT1pGuHGsIZjzC7T8QodcnVqt/Dy0ckzbluY
SLLtdxNMXt2iLdo0gdweIncGNOi7+NoxdL7c9HU2zmQ1ghqhsvsVwK57a8Y9fHAi
oA5EguDZlpgzV43USGdNpPYI9LjaUArwLnyUXiuR7MSB3/HbIED4xG5iWTRaeAvN
coVg5ZQ95EZBys/ia5Ix1WgAWB+fAagjVauukOHXb9ELGaUlhOSpFr9Gvl10NXyZ
LQ5ArGVFjmUbmMrA5TRmNj+zTHmhWDwEmrytccH9kXfqx0uD9bJEp5lNkh/FeWS9
J2NviIY5NB7yQNIkxOWZpgti8X/EkumdSKJxVzreBpGLedoDFblCGKsSzQQuM6SI
67LT1oK+UGOJ3Pj1g+VQOPafK8EWUvX1PGZdZ/qnuAr8uQm04QcKbC4OPxIw31Kc
CmDbc8HIcfS6nJeUrvdxLLNYTWEk6139vcCR1W/kyrn4iRBvJ3J6c5QTDWtemvXD
Iml7Jc8JBcFCJQL1Se9VAjOD29uDB4G4DNMdeEuCONLTrzafqdpGIiGlSEftozOn
pIv3xlugVh1qCACNIrjTN3QMwS0tsqAx/WcgGVN3RoJ5OYVVNh11qjm0vkfNLn3I
kh29oAl0hlvZ05gujz++bJvO9uyqj0Ot8AD+wdtc+zNyc/dbsVfWB2eQzwFLwiCZ
I7Ik+5w5Vz8k1hU6wTdg6edwZckBOXTr7Epe6keGKCgd53vHrMPYVLgDNq6fpzoe
qIWXECgmkWPLQs+6hwVfquD3rTNlvEY3dbbX4gHrcb4Z5MJWGl27+ZMdT0K3t8W9
5Gtn/TQuZN7kfBUvdb67oN00VI6pDrEY6tI3CkkGQEPVZAK4ArTX2tAjFxNNAhJW
EXRPFGAdhEncYvQhRl6c/j2bRCom3V2osyj1yIsSm+ga8PHJR7Lg2AMk3uCfGlO5
QdHDasIoFcvk9QdWsAqdVZg28CcpfOJ+eJESrdTkp70BqxfH477giv/T0h9KXuOs
TwhKmsYoz5+uo4dMa/zYTD1mCWOr3LJ9Z8A19q5xW6ZJe9WjXBZTunO9H4gAGRiV
/nVlxsLeKEgLX+mbbYtpqgSVfvmg/FrSH3UWDkFVsxB7LMa1pogIOcqrK7GVw+As
pbm0/xjAFe70XU1bfEQVQ/QkPcDQRC9WgfjFHzk4uvYaPEA5PHihxzzTh29Pf5up
sdcGv9zxJGvIYMwELVhvr9dS0kQkqMuCn65qYilmZC++rPFkTpnetVvajeaFi/VL
ngPpDtjQu01sD3XQoCwFpD8A9gPXMtH6V20Vv5DMLZIfLSkbQVNZCtHwytx1OJJC
JPfyFOyKYFiTViUDHTlMlVuzTcHhM1kST5g4XQS1eneELJf2dlLeh9dwvcQYpKoW
SAkUSyVbyjxKBg6CDr2ap8L2gugXBpUClWezaFHBR104pnkQfImaN5uyMmZqTsYx
a3wRPSVJr9lWMxG/+VhlHaaXUbr7bFftDqtm5nPTryrGLiyhbhWaiRIGAT1iZC9R
X0oQ3peUVNkuvEQ/nWi286Qr+2No3klMyu/2GQvuyoKwH4+4btq8ts1g4rya7yH+
gounLKX2hA2IvD9YzBc+xY7LlsS1ETAauVLKhBDlvgGddezOZ0GCx5gPPXb8GZDS
wYuKjQ0nIQUFSLsiOV+Qr8C8otn4/nsGgleWbMhhQC+MzAsMw23/AlijDAicgsDP
v8GBtmvoxXNaNczbGU4ZR0ktcXukd6hb8RWWLJUXaTx1y0/IaX4x3Nc9uF+3Cd9I
DGAE3zz6ccgRlEi7SNbfpTHmB9HiU9b7HM1n8oVSTeT6ck+B0MG5ZeZaWTBZdVoX
8hqmupqgFxDWs9/5Wl+7kPqzIgBt8tQ8NKvGY3hfbXY1D5k0FdDqJojc4KhFV+BB
XVYn9fBYwj3yjT/Sl3Ac3ccxHGXfzJz7Za11cyWQFpC3fKikNQkfzupFGO5h+ICM
frmzYV+35yJMkJ9f1wI2wP+5pdwOi1MRf+Rij0JYRGTbcq1w0AxE2nIY0Ltr4epq
J6QBd/+A/TMhIttDGmF/jR81Hsxyaiwt4Rrc7HyY9dO/WiRSBV2UAYM7Nylj3/Xy
KQi2+hCDy43Ll3p2h1OxHPQYQPnGdWTNWHlBrEhSqOJY9ve4I7YAH3/B1Zz/rwHf
Y1Kk5K1cZCnU8UVpzBwRXOgDKMFRzwOkzeu97VmcyZoza9puKrnMyzP8pjQ/x43j
ZeGADJTSp1gTbQ2ieroNonfmSu+6tEvqg83lweRVvCCFXDVfpgd5LYH4ETKXH5Yc
ynIY1FJFXmxoMUnJswXmPSIIFmRMpQ1s4cQ5dLlmN4Zl2l+eKEt3mp5tep87jiUq
EX9i4UYg/IxQxb8JBGR27LMWt2u8a+V2jKoQHRqdKnUJ5wVRANxf5J1SQ7QZpe5W
zES/657KdSELSArFNMlMIwQFHYLfPRnybClGGAckT7SB1dUEulz90uVrNCfupEwN
RjgreywJQuCvY5ycrY1DHm0COvydfdK0+LjbyhBkZnkvInCCYhtP/GNy8/6B5BGh
ux/xhChD6CHOsfdYpZ9OosWlWLIZI5ECHdXEFcfSXtJ5VU6xxaYgP7EdtCCS6Nwy
HDzJCSRZVPBe1x+kLwMdjTcoLLYzqqzuM+JHxfUyfs7SwHkdm3lgQZ+ry0APDoCh
oXRtZe431ASALD8meg+RJDDhYS9nMqcrq5eFmV5Vp2wtixjf57OApf375ce2+ndx
UmVZdQLmVBDB5TWzo8YPU2tWaMs1n3wPf+qki2hhGZ3CP7OAGKIbejGz2jw7BaZi
3T80DkcPX5cHvMvPiLVDCKhXWCcmiFkZk8gQFS0zmCWQF6RA7f6y95Zi8OgWxYj8
4+LAmA5pbyy/JWfI4otAxhQoBZSDEuyT7V4euqTiFqRJiG1nQPZOk5Z6OWtviPlO
WkdX34KuxQzux1Rpmey4yBUKLtIORevQ1Q1onxmmctgjFV49kbbOfhG/1aVQSpu0
vLHWMxZ26o/mkh5qJhzrl+HvuL7wRXyYxyq72xiMn34kdhsSInmXr7xluOk0D9UR
NB8lXNshGLWENlVLEhykocmi3En5xaTkBXgi8omTv0LQ+R5QZtTJq7FJ5cAjc0ga
ngwMHbsSQBtmCCGvmCh3NjpEqgjR+Yz+p01hpseB/6Orq4xG5qASse8cBnEfCps9
jvn8LGINWMMtDL6IAiX3M/J+o42ZVcauFgEidPv/kd7S27IbEZj5WoaMI2/NkoKg
zyZSyRequ6YTo7RCK8L/qDIQwIZlQjpM1hzuL9VJRrNbR/UbZbU0CSPMkjxFJiR8
8rZJBMF2ao/LAmZgmgxi/g2Jk9Vpqxia9OBycZuiCDiyNi2nvwkR7WLKMKZq72Ew
4cVra8vCehCvXLhBY+eAzR2cZMdo5S/wWmrWmB2thNolyKwdehzyJYDG+THBB352
oHLNJFCg5V+lTpFWk0yaenn+dURQ2aEde8dVjb/vmSPIf8CivSVw5Ot6/0eVvM4r
VzHRGPq8uuMzAdwzt8LTE3mst8ya52BHzfMV4CMKRkzleNMWf3/mimLpf3cubbK6
2hKDbw2m4hokCca52bZjmzppu8xZUxqvJ5l8s7ga9XnZ+U28EpeVw0zCMPGr6PKj
6pwRS+swyrLdVfVuz30P+o1YFcfWHA1DLSfD1ZlP5NbbguTeLdlgfo6gS2nqfaLO
d6KxsXqdt16GVudpzhXQPl3PQLqVw2xiFYMxv6dVceYKbARLlEqYFtboou5DO965
wuFbCHTod3mRpofRoybbWh8Ia+l3ao8FEfx06WBxhZkSFxXO+VFotznoQGoK2inm
4Z4kRukm8W0zCU0p5KslLHnUWN1BB68BCqNtC9VgXt2etN18BVz+HUwdCP6hVCoL
awwC0Y2doUQ4yhDJzkQTw3Tqg/zEcW3afk1dUX+9O/IU5sKAJVsfWFZ3QHXd26pN
r9XoYyS0/OdFVtIISavxm0GMrXvJ22Wwd5Q3L55xa5XuoEoYkfUp5pTCJxZdOcol
pruoDJTMCoB6lMHQXOYgtxIvUrk+SN2tX4aE4cxrkCyetD8JrjKKfTv7SpiSgSGL
L5tlW0qTq9R8zrDBXTpJNEF2N+X8I/rU8kpyNEMNZVVFh28siVRsvfZcsiMrJRyf
MV0UObCnAF7u4j0PkMvoclcXX/c66DUojngA4RnvpqcEk2UTYiNQ+Zi4y6HmeZvp
gquB+H7pM8U4wd4/Cb6hTa2cVDF1IYVYbq0+bzP3mEIFRI5GvNOlMAgMX1FsDjdZ
FJCFqWRo6sL49bL81ICVGzPmuMPgmWafbxb9RCdz8cR4aQN6hUmWwlJdeBpp8ys3
X9Lh1AtydsfyxyktbEJjOTR4uLrjy46KHSrjHi9N3aB5ui99Kx5WgRSik0WbT/Z8
x3LTlMzdjcbK/YSLopUARHopzO7cH6w80ni17SJBYl47KS6XTqn4Citn8sKtuDbd
ffyJHXeXyNJhaxnAq7vv3QyegrlbQg1UxABKUX8dSmr2EObxNAciEFN74pyqwtze
W7gNWm4KfLHnzGCR8v4iz2BU3fRb8+xvtjKzguZPThHgIE/n+ryxtr7MipZ5aEZU
t6fJQFioTaAJ1qbsYiJeTguW2MXTfciS5LWfe89Du0Y816ZpVMuDyTOymQG5zaal
ceyweHAnsR3Q11lPXrQzb4Xg/BZ1/RAZBphPo/jeBABUEbYt9tecs8bBFpNvyv2a
P5G+3jbPMLQq6Hn/DpIIqYFlHdxKJRcrjM2fyayGSyVk749pgQjF4Cd2K/zCiUai
lijRqJHf8bvCvBpkEMc3ob3UIe1F5f6noUQxKvI3fU7PEoT6Fj5LPe9+Vwyq2uLF
rBlqmfgnbYCN57q5q5y+Nyg4W7CvkMC8FBJTYmB8StM2eWB+IDzoWmXfLS1ot/Wp
3f1nxILTzAbfnpKBYpIm4pGsfI0M2tvGxCuR1YG59DoAkyPMy7h3hwAkr7vGiLNV
mVIGle/t5PGis3WYAsYhV43/xJ7RjxJKCTazXpDHTClQ8UNUBCJyE0c3UZh/atfF
fMb3PjvZAdL1Ycu8JviYrexz6cm5kpkxgcCOiS4VnesMSJz9kTH1NctZDS3yxgUO
TRRv/swOJgLmx0qaBzX4o8xP/Hj4KrGA4t+sRGpOAO5c1Kmorau5dH0zrT6AUcVN
JLzwcVuHi5ukqC1tVKYC87iqdeVgiLVxWwsKfoaQGpOX+P4c2Abxl8afBoY2KUtJ
RwdvhD35m5tROwGp5afC8onjFQ2yvWMFJVsk/cPamDHSANhl+KVrkXYB0MYTLUmv
n2tmzz3PiSCaqNc292EMmvEcSoNa2dx7nY0tnlcHMWqjhp9bIlvH1yNdnJ9u3cXZ
kk1JePWXhF2moS645tOPENlvwAfvr/6V/FiSJr2K42rmAJC4meVMUgVAIO4wZfcg
Z0CirvBsNReA97Iff6Goe72S5vWvc3Fiarm1XMdjnwjCXuG7fczhlGzyYOueYcxf
H66eNVXi8VjYkLAx854hQJlYLiYnztIHakBfXBGgyRJ65nvLYiI1NT1hJTXeYXMI
CZPXejrgaZPur6JI6LjQ3N3cQ2iRe2GbinVvo+E5NyxxGcvOX2ljP+otKoB1BJh3
KRoc1w6w/CVaUQ10XNGEcuVyd2DKAd8ZNLCxlxm0i1DqAfjrALXY0wQu9FzgjF1h
+NjJUXIkKiByY147qkY1YkRZI8QMfpJLBWfrmEP6RbG1n/lvoTnNoVbxZJGsDPD9
OYzg+5IBT3fsCZP5AU0qArjDbE533iTaO6dH4pmx+6GEEjfAqdtoNXwAj3NHMy/Z
JvhcHr5wSl5a9+rfvGAhSZ9Lwv9Q/o9S/RgA9Qze8viUwcUsScx5MjW868jkrbT2
VhmobmZ6JgMFQvaPbBm0psK1IDoqCj4CBKGKWV01CZAaCpsahXfCe04YRAW4eHX4
mL4R0PyE3tw730zNfv4Follo5TWPajc7Z9o17Nbm5iuJ589RVvVRorm9xHacEzS9
AmZceLUKyT4kNHVdUgLhgxKq0aJ1THQmSOesmei3rT2LHDpAdZfaqvThBrOvNAVn
y+GHWJ3NsNJVGKm8V5X2ZmpA7HHDoVwoUa9cmxjywpg1DTuTx5li6dBjV5Pz4EK/
BuUeWl+976z0bwZBG/7n0Oj7GiT4QAZ9jwbgnUF8u8p8SjmurivWVVDMiOuiiidG
ptrmT/A4yYYj9S2CtnXzPbv+svJGsznZnCpQdfpTSF4TpnLsi7oD9CZHR46FyoKF
On3gef3TjRUcPOcUr8c7qgDnMAZ5n8+4oze7Qnw07Avt2H1Szdy/2sE/+np46GkX
qAmdpszwt4qcsVJ2P27ZFzDZMgz3stRWUe7QlVyyV2jWwSnldLS8XQaWduXDXtXT
hiYJgg9ffG6+YLzEiMUlqrsRGeGeYwtvCdq2wqgsArlR7vVkRJQ/1j6kwWZITRst
xzanGqbmO7nOb4RhZ7uDSutV7DxvbpjtlKnc9QVNSy3B9iW0z74k/dWZgIp/14BT
pDg/QrVUTLi6xKYiB3WcdOSHFX85aZRdrhkd2n7W/khBP1DWhEffb+XEg4VMMqLv
wvYvOfPOTX0Q8LO0FDJUZzxOA+AwbM9jRGArB/C5b5z8e5IlFJOKkdUFf6vMXhM0
AD4kGLutX6MVQXnAQPJfoSK5M/OhU4UIQjc4Ud0dYuGtvL6GfFGBg51m2VKQO2E+
sPKiym3o+Pi2lLRsEANPY1yyWcujOunH4whKMNFGD8dzv1EtIPRWh8OEdWdJF8xd
EMQH7Ij8nW68oxVdVI6IV1lxOm1esEO9f4pnbIYz4sJqJGZI3LjWvYvzYnfiHVFk
wiAiOzfcxihZsiuMa6i//rP7sPSDcs08NdPuHr8HyLgQR3KnrBLY6sjjpf73ECim
XPkdF6/8js9VyGdMVERlIdP4i539mPjrehsDp7jD0GifyCSMbAE3qkLoLE/lcqgF
oQtQ0Fq6O0T0NIMKxAh0eR7sEuUGhqiop2VZlko10Wov79vKZUzv9241KC/WuD+2
R3X8zAI4rGfvWkKevPjeOOeDAVvreLyeY1yUAxVScl99gNVIX7afL13yRfangCZc
ljNFOWSYy7BzeFrwicugNnQ0zwdgXk0z92fSUHAztDzvIb4MpLAsIviZPINrgx7V
v0BvXUaa1tKz1+2R3CiYCti5sDhYY7YXqaTEi8O2ixY7RXDF7ZVIu83W26sya+CI
5qNmv6JF6Hv0w68XgF9mbz5CHqlhWmcIIhvz3Ti23tlPTiI3QOp4oagQwd0+DEwK
0PqOlpkiSYrt1huCWRozonnLW8QV9OGFdZ2QElPA6i2AEjnNdhRWCq6eutyCPoAO
OZKFFM6UCs3c1a2Okfyz+QChEm5mkRI+QWdm3UPEab/EKspqBenbaIbY5iKYKyJf
qqevcunnBFmqCkD+JUQEO1fhqOFHMJp3k3XlP0CBzEedrj5rPzsK22qspnI5ybDl
qUjoGvT01OfhR8HOa83KJ4dG+MniUg0QREXeQgBCSKFvms7REY85B8Wa/KWLqS3/
cL4PQFXAI6I/pbis3UoV6BUV0HEBQ1h23rmWX+LYudFmgWOSabh88busrjIH7eW5
axroQwESHD2M6NBbfydFT/UMf2PU67kTS9t7FrKzQbDRLiA9scOsjc2TpfW8ayIK
2YMy+KALqm49M3VS5R0OvmBhbtbmc8KJDZCVb4EmFvB8gA9Q++Z30+oj97FFhU6m
Ur5KlIuTpdd2bnGxqakbYI0uzRcMczFr5rDyYbnmllqwu6KdAFAZ8NhLwt7YncX9
MgvNAay2LA8UAOM48qK/qdfifoRXvPbAEN73b2eNu782avcl7QWtVpwQBhKvy3sw
2qun70ERS3qxF9L9yd+IArcBcNCQ2KkD/Ka3UAV7auRl70kQRRV61BBUV4kZY7mO
WYxvHsmnptmxlPJ8v2VdQohHYe+SAE+0fUsVJ9v3ag05z5+OJusQXfayiHHWDVXP
pG9jnvRGmXN0uSjDtRKumwNQFT+j9i5U9PP755b0az/g64zYK5tR8V0g0rIbzF5B
cG0yfVA4WxVd+OAmV5kP/RDunF9qoInmaf3DKDObZXBpSbH9VinjzYAf/nRDkneD
L34oqkSdg90Z7/P1XVICoS/dexUy9cFGkwRR7+L43xr4bTQnW9y8e7/uwHURWHMQ
Lt0Gj4r9HpBFnnNboxX2+0tEylXH96/fzD4GuL0AMb295vcNXXWTV9ZfCP+eP9VH
Au0wY3duaIx8UTFF89HA3lQvDaBynntI283OI9ySb3mum50ECA2JU4iY7UUfMR6R
PoeVbfeHy88YfAoBKZWH5SSDyTvxWZmQzG9DqLTgVujm2daLJbNcLTC8IDobjITD
CRdnk/uegFhR8yiLHUYXWcT+a1M9nWG4BlBi9LHrj+zvsFCON7taSP6vUzd/zOjI
CUfjSlao2NN3er+LHVGMdmNZn5rvnlE1vcz2l8y9Ferlzvf2Z2PLn5F504eVST+S
aYPCXVC95ZoYhporLhuCP8rIRj5gG+y+MBqd+/0sC+wiKfZn3gHDoFpX92a4Mtn2
HBuNSUUTyyUdf5SQH1yymjAQNhpUs79miHJpnHkI1AL5KV0pGSj4qF8gSBbd3+1I
N0nd9Vtmf2stKpoMBiSMcf9c3/4zd4G5slkPzUtdRUzpVcEfb8dwxQkj0BWbZ+z4
prARGTVlfIMNDkc/uXHTRElPP8JNI9whWPCrqxZ8MuPAucCfi63FU+gpqhuxZI9m
v1KtltuFZnqkVRLC0aT+x1bgvBcigjEzANlHthidx7kGeNcKoYgffNtylQly+06k
xFuz0IQnkz6W0JU4lx8xy2nMNJIw2H/hz5zRMTgBy+m+Ix6wUXGZbFxPe5yZWxUw
a++qqUKQ0q8eDP+l+VHqMkid7DAiY+6d16a8+XPX0zqf377v+kF3Okb0rNQWBOJy
YpZT8uqrLBDkHN8S2LiJEB1ZDuyLF3CsFM0jRs571G+KLk6lgFqX97gz9GXPS/IM
Ut0fmrBbgcN8SgNkihiI75mhtX8BYx1StI4xHTlAfyVH17APA3Ekhb8OIlXEUye+
rKjXG9uXW0X9FzWs3fNspD/sVWJqiO8YYijL2pDL6cc/E2pH8SsC42tbgjrQzRUb
Ns/3UE3mXfmMsf9lddUVgJm0U1LEML9NhAu3H24JqmKDUcQkesqWk3bQ24KBZ8Aw
qSFPYUO5f03HMm02OkjeDL5jzqmRUWeaEsdJfH+cs7KWz0ouqtcEnBHU4reGSSm3
NbO9yoaPdhbFnphroahfvnj0MRfepsEr4nSaODa5X2WDnV8UXKCa6J9WXonxHwoE
eBkUvn7CqeLjxMRGFFLoVj0ba+M2BdJqCTeDGhnhNRkFuMyEcsZ2f7anWCvMFqHi
XanYpfnbXZRfdPkgrce7gXYlaiIw+AuajMWJsDgtlWP4q7dU2V4MJuwPvE9qc2Jv
BKLWtTdDesZ+orvFNNMTO978vhuIuOsVcUWDfhDIVRVhUz6VvYdDijRIM1F3RoUG
26I+UFVmhv0d568wgYW3PXOFn0szt0F6Rteu7FQIjNWAsmig6+rvgt+cRkole8lB
GGyLp6FPq2wtbYbXx6olDVhe22TxZW4/Z604zjH4lX90FzhK1Sm+jQ88+93Z5Wlg
DDpLkfJvXraJjaIg89FNMkljMCnC/tNBg7dRs45HbDjP/0OtDHSr3WLR5dJJTLwA
UxLTl0tOalNi5n8hPHhZ8aN1pWNcJJRP2XgkCtj8c5zJoGGIQDpCoazGL4x9nSS6
I95A3M1UjvdzZ8d8tGeAIhM9SWfsUULofDa6CgIcv4EYyfyTRzo09MNoZvKWoZdI
CnY6FOeWvvHDd6ttxBYsYWUjtDWW7bbZqKASc0x8s5aVa1XZ6W4bq/hBHBbmftW8
KR7QeJ+lj0pTdGz2Oi2dw/Z3DDXNxRwhcld6rhBOxn2J6UDVUzUqxgDR9fMmxpGG
4Of6Py0wXfrGsC2NeUtGAeU0P7qZJuqIv5XeXjWMv9Ptcvo9gfUY0vZ/d/GbTvLz
j6cg2TJJJi+WpzqFcMgjXK5wmmkfqKyGWOSgXSxaU1tCmOGqLpdgXFjQtF8JjbuC
TUm8BrjaaKtaxhL4U61o30qajkZseTp5Q81pDFSqGoZ+rXuW2o4AjGzrsJycDn/T
oTaJyMWNwA+e59v14T+ZjBuyhag5m7gybmJKo00oyLw9Dw3Qxf2d1SraPTFD8y0v
MVmNywaAvcmBS2HCcBTAfM8nwnkS7WNzK4yCM8Q9eCmvALgxiJxDwCaQrLiKYpHc
FpWjWXeYCcKc8Q5jIBEOtPrnU0PjEyfNs9WhAgQ5O9y3Gk/eBNlT5A8uf2yjsNgS
zMFGySWmVqsJgoZcm75E/gped9Kzd15PofTBIjkq7CuUHpOPjFZWybcqPreBBA5c
VmnZvC8ZB/N/qm8KUGzHvV6IfvqNubX3I01UnCzAGbPxv04vGIFPUcQ7IO7U6TZk
ws42ZrR3dliPR2vYvnhCEIzvNb1UabI2C7wzQliQMA3rz9O58lOpm1uAsxkVUA8U
EHff/KhshboFSDiICN9SsjZyFEPW0k2ByULordmph/cI3v+DK9NVSvwMFPpJMeDZ
eYL2weuFD+MbphfleFxgodVQ1UWOuNtmVMG6JocQfaSE0KbAO7rfOBGPzWDI9JXt
/HfudCGaN+NeyFgDpeMFzzvfmm4C2X7JLBBuVzCpOMm8Sp2Yd6mwIZq9UMBCku89
B8ifPHYuaaVKoCwU5fBLODvqOL26BTQHGXdfRa4B/J2oLZoovB9IzoJwrm7tua1Y
7LykbQqrgFd568OU/WALz13x5yrK5mWXUQeEfgQyjsKZdYVVOSlKP/fXKFdnG/tI
xet7WIi/ql2FOtJvIdHQZLIVKfsjsamFjHtHVQE9YI01o4DIF5PaYIspEZ90YJVh
Q2Ev8bQZyb1meMv734ee4Q79ZWfzj4C9k2vOLBpCBViMYJHvMOj50jkyU7plAGN4
cAa/Aw03O0F11IOA61rUVfjpiohGqkLP624ih7NESXyNTg8C/21lbv1irlfgOYvX
+yLwPn3nmP0GFQfnofO4NIWxT128RY7/fugnxHayq8gCWE4WiisqSDV/m7AiLapG
wQhLL2B2llzsAKfNQ4aBJoG4XbKXF8lN0f8FkvAoFqUSV5wluxpGMFDO8l8nVj36
aWOahrUg3WVYdZA8smxPob5xiJq+9f07l2NJ2AZjMlg91z2EV1wUK2mn9dnNddJn
gjXZ/dHlidGBjEpBgq7nWJUA1/SqCfZf65UKxD+dLOsl1iBWBEMUYUkWQjR6+fkt
lCltbyoQft19KyVzoFPRjeOYWuZHWZzf8pTJa45mlLX9/iv8ylOeVO7ZxikuxH3x
CTglo+j0Q2USW0cBlP9g4TQe41upokTRtg5BrZ4hAXmm5UCtSQjgqHj7SYzCJvh7
qQLlbtQpS96bacCVdzAj5alBFy45Xrwi/qUkzqEcI/aHVsg/r/pxC/QhcYY6XaKL
EPBWeFwGLavrsm6lHR4pTGHh2Iu2AQD149Ks+gEXH1SLyRchjuYUJPWT3gPOA4mx
C3enOZ3CBZdQ8WhOModi8B4UJIofBGTsdGwVRctCWunYRXRl4v+qH9fh39xhcIr1
q3JovuWbM2o8m5bdNXvsDd1CJRxwevLmYy6AqWlaeNADV8bjv8mqu36m1XlRlddY
WDVDRmCdd8GfZA9BXyqor66NAf576PI/N8cz+Rudbikw8PgUL1KOkAImWRg62tyc
9h0qEdg9loaq40c5n12qwaDQsYmfZUqO288/MDip8Jb6i9imCA6cb7TdyiZA9sId
5l3SpUOuQnitypT/tPpphG86DrmF2yCz4WL0u0uBrwbEIn3eqDoMdpdqkftW06nb
ty3LIIh1xewlcUlPI76Tm6nNz/YJY88NdpXBAkDWwEX9qCfySt6zit+SmweBBSjz
L8ALK1C4eFL2VuopF72gg61SwQqx0i0/W3WPswDqnjsxKjbZa8FZqADdl8VYs1i9
gtiPgbGTuiV4BDrexo2E7h6nOGoKK9wWooFH8PksjbeUqjRBogVC3OtskqhG1368
druEMi2CZM+PgUpw5tJOIvknPg4NCwe5Zx01kOl0+0RkiUTk5mtbLtend2HuNkwz
5rVVyuUKmmSJB/tKs8C6KWuctDJy6oRXKX1/Bb9On625eLohrSi5kgpJ9v2/iesI
uRs8GGet4HtpN7osF7IUMh9ae2w4mBoe087t5rDGOzryT+piKivooc+rno0L6TEz
vTNXDe6szZBLnoqef2LN3NW0Bgtl4+jlQkpSZZWWuBZci1p7O5OmzYb7HNcvPCWK
fIjGdpRDFfpEj4Nu/Z8VgkBvL2/OMt8qy8fOOnteeYvkeh6N8iHYiuVhagSHqw8m
/VqE8tFYGBU1u+4oB2KfEqFIbYvJJPT+hRPxd1bRvEYNVBudVndAtmQD0sSWxIqe
OS+auLpM5INnvdnRifIfZQPLflHtwLhvKhItjMVhNjNveRsIF7BEIIOrPbKl15NO
ULE75mAswppAhOVNsi1WdQ0eOAIe7HObO6Z6BxlxXhUFMXo2hAu4MwDjt/OI8DOi
M82aDhEA74KSS48QTsXO5T4fpbpB98qRBmRRQb0jAwLOtkHM7rQ9npiZiD5VrCcF
Yn++o0Lw6tUQEa34/GG1wU92uTNtoJ2QztBRBiBMEjaIQQzNtv/8S+ZueFODIimW
gIysc5Ulq7jocMHc9pwdRD0MdQYTa9Hlv38J/gvAkMBTdcwwVrqkkXKd/lmslr1+
5hZFle4NvxfJkycwTNzVwptpk2SV5gabUVMjDyuc4y9EHfJWlvL2XqaNt/7XOTLu
bhgnEHhRS+2kU5f436G7y9w/VNc/Ctkac21vV6Ih55nt2UGICUMbFW143GXP6sAz
m2bhgXxKdhe7JNJvuBlhrnwRg0FREun52+0xmKvxGtepJQjwMEgHsuK4uoCMKnne
VkFC4Xjob3MYlda6z/GYnaVvOO91W2rAWaNVCnV+RgKTvPXUzjba+FafF6yGL5Ii
T5XMMV2VQqJUjePzJezTQXEM7ZUFXvq/kj7vbwm/w7ISVws2lXIA5sA5UKkf6W3s
33UHo1Oj+bsyUMgBEm0m56s/ypAvM0dXAFRcdCE4uNywoEn2T8yr8NF4hn5ClP0b
ClUhAqPWDXkfb7qPIBAZC3GYaAZrfnmGJu8kZhRE/5y3OKQP4mbPVDAZ3wfi1kSL
sB4ryf9z5frHHzlRh89Ao4Q1sHATf77QoPJaIU/Ha9kvI9OkBMVbfywxO6r/i5RX
nQWYZP0N1tpBCwdz0DYds7tmLbS64KcO5HxEHVYxdnCCXt5qv3chjRt7G8eMDV4f
G5wYlmkIPks3uKDhdZ1ZT4OEAANOgGIkoB8oirMLt/jdRTf+uUXcT6DrneZgTqls
Xm+zrVdvvH1O7JsdxDvw7j4vDDNOsGV9z8Nodj6H0G62iKkZmjVTFGumfeEMixgA
FX1tEpM3UYz4n9fSEz3MpO1uW5hoJyl6ZWWCx1sXe1fNHAZksjcfov4Bq+wvu1zu
D02Wx2foyrXg7u+AbOJkmJtCJYG2mhgANSawlu4UZmoLGqjkgyv94OY9W4rigDl6
NFWbetXDVTr3j0g+ldff1V+e8zagbbGgc4MZ9U0r5wM4job0FdUzoN3GBIDnThOm
I3CqFzGNxm2llCJx3BOgcBPIXP+GoxKgJQT2B4ut942d64hC6Wb1em5DQlT1MTjs
xEPUuo+0tWs6gDajjS8WQDersc6Uf0/W++i+q4Dp5dY=
//pragma protect end_data_block
//pragma protect digest_block
hXe2p+GJOH/i41O3HHQOReUR2nU=
//pragma protect end_digest_block
//pragma protect end_protected
