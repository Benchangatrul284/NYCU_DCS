//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
ZZFX9RUT1cZ6xKSSNXzQ6bnhVz+5A4+2t6hcR8gGVAfom2OfVnD8CVuhDyGBDK1Z
4HRRkCELwZrypf5y+A2Ioxw7Fp/QsxePoNl7mM+zgzUD16BDithmwXO6TgZthgM3
hNhLToQ7FJHaX4Rf2s+FfzW0PL/jAlcAFvaGD9d/PEHlYHmr13koPYe6L6I4tkWG
j10fcg88hnqhVha9VjzsRoPD+n985Gu1SekHoMVLb7YRvMRKF8AIz49nw3lCzHZ6
4acQjBxztsNjdcNl0u5/Mz6FUwCqS47KybH6LM4wXumvdQIMiKTsl/vxIPUyCjt3
FJZBSzXofGPsfaXyn0TSuQ==
//pragma protect end_key_block
//pragma protect digest_block
ZG1O9703fk6mQqqnNmdkppUmKPY=
//pragma protect end_digest_block
//pragma protect data_block
K1Wi7k5/ci15bCoJ5QrvZE1rCXUWTKkCa4RRfxafa7U03RLpTNJ+HF+naUdLu3kk
t2GKPXp+avDeCpgnB6M8hWPk32bbMy41knV60iaA1X+TXZwYjHSR7gp3dkmdHvUi
KjHPpUoMLk9dDHti43O7dixxNWKW8yJpF11PDULVJKnTsVNzKM9Qk7l5LuIPVkka
eVcM7nyR3nNYhr+L/Xr2I24lGb84WqP6gfcImGvS/+ykB5aUrGjylTDLZ/rNcHui
z0+ReDIg15Spf/zmETaTpgseJFiP7clDSoYm6xPGboXqN3Z9/Kwipi6xdHTyQVyE
qP7GTgU7WRfFBs4cnZJTvTYXrpR277X6wkbVUtyBsTOZE8ORz5Fhuq8wp1a48IMc
YaV7QZltWhBy1HZkSAlnx9Z6uhztuAJ+MZ97zBdRLTmfCHJcJkhj7x8JXv23bndf
ECrwz6zva9I0YVmCK2UoQeOv/PfpDcYMnoUMuTLpacXDDmRY5MXW5AfCEfqegiFY
XzyRLebdXWbnIZWpzA+zaEwyHTVLyBAl5wG9rgZ3IKBOVavFpIX8F9m/79i+whC8
cwiiEw0bF25TY5oGiyhN7Qvo63m6j/Y3vB2gC5IiJlyJP8B59ZD/CiBJpMVOYr1x
MI3+oHvArwCRcGJKAuZLmmjCs8aVUcBhnM1QgrmbQinOjNphO5/KamaU9fczcxoq
3kG3yWgKf9tWGOGV6da6pqr6rqOiEYVWyGQu/uH9HEXDF/LPSGZoPk+oo2Bg2Tpn
j1QDF/a/YcySS5VSXJmAvOo/zFSu26gMhYyQiZT3mewJkuWUuEjrnzyjTondy2KP
pBOuwMRz+zV20SNY1rH9DP/jYK3F6uwnm25cOn/Y6uCzZ0XkLq55br2Es2Kkr3GO
aepQZmixgLE1AjCHhL0qcMjI2NnoQAFecuYvRZSf5rwFhuX3qJTMGTcIIkfKNK5W
nkoY0/qGF9yj5iPNbMmxdPitRu17tlThRbkCVA+oH0XPFHtK16vGeAq/DeoxqfoU
CiHJrPHKXDvte60uzw6OM5ZJki0HK+hSB+cCjvxpm1leRBbmYWb3zFiMMNBawsWb
v4mqt3eP3KMC1+VQqwybkugIA/pUREQsUDqCkbdp+sZQ3uABuhmCuVkZ2c+bufEZ
klvRkWFALxVbJpBznOsYGehnSYEG6pRyJyC0cX2WeRqtX7ZA7ecjWtmYKiVtTlmd
Q/BC25toEhwU9oxamV3sRvueJ/nCa8FmjXAzbqUIkPtYGuFBZzXQoMQgB5hIlInq
8dZAJOCIvfNKLpYYwMt6Q+6PAMHeqTC1HD6lsLJ9j+Q+7n/e9UmQvKQwcOFXZaEO
Aw4GTz0wWmls4owFf7+EKMFxNzleY6HDB9Jdn/6EYp186MRRfxdEEdEESb2VhnkF
+OV/cB6hWwXh2ZL8gybbQG4cZhP4EKnizGx7b3p0gybB/aWAfbRHyhYOtDu75Qrs
MRXAsZbZlEuF9HeCDzpdRAmF7jsjghxxTtjkuurhK0OPk/NgD/6v+cCPIb3FNL5d
QsTtTvtADRugTNIk2YD3MA4zExZt9FsKjODiJuF1sNHvWN8hdNQQ4YB8hxECAsHm
t402Aov9JBpEwzc/DONr2LnrhEtOCLZqtahWaP8t7SgxeZSGTdUvEF6jPHxMZjv5
7cZnHFGz1umxHSqjQDB7/jpXDPB/nzFT7l2PkXo/dAwiOrACvsvx0DPaHCAQaplv
Zh/k+i7nMTHtkx6MSA4ydfECC/Bh80HFCHDpQOnC0XkFcjbuiJ/klGtP0wFciLQF
W152A478wEMtSe2Wzp9Cmbq2g4WLY9LeeCqBLWtHt5z5ulew/86Gg9jtEZIoCfi8
7DUXc7WFwb4qbJxh5TF02kuPKOshucdrExCy6lIXs5JE3c4zhBDurMMd+jYjVKvL
S63seDrW2xgDrzhBs9HVEvK4xUXifIN7tzNocSBe1mc0XziImK2w8aaw9tJVt3HE
pLLDV53U9PRZ2ETy2CauSd2KASxZcAvb+dlzLlq73huzeavcnsx+V0nIOQoZce03
/wUL+1AZ9+GH+Lh9KoUnW2HtKblbUeh0wnQd/bNizKR4hQAWMTxmQW1Xj6OMhYCD
eVUUwpAAHhE5ZztEZzi/8wy7x4eGJd0D3uW4Pg0tOXmDBnqVUXoG9RUmQoqGWTrh
7hsLE1IWH66t8ATu7m6s6WsqayXI7+qFl0M5TqfBn61nx5+tjcgKdzcTNkmldJxS
kbP65cPFMe2x28sEupD50CMNUcE8PsSpUQUTgup+LgadT338Mku57hG3Waq4zK9f
GOlmDLXF0794MZngBG0Mvev5qTOBdIjdNzFi8G0TGzAySRbaERyEP9rQQT2HrvHv
DmaYJyKomT6Xiy/dFspBJbBJGC+nDXgqLHrGz6RpdON0+XOOW8OUEr1oxzzrg8xM
dfs1l7vR3RxdolgYMKYf7hK9dB23527OcTgEl+NAin12HNBQ3Pbw2EyBeH5raYCw
QJvi2AFrtdT3Jh7YnDZMz7IpjaB1opSO741So94VRyVyGPwWp/+2WFi3TQf2gqAy
5VciCQZyPny6pIqFELZNjlU4OjnoN4uLX4fPEFlgUc2/KX7/Vs0nNpCxjuEsfu6m
cUcgCEsgrsmhweUZtcU1QfG8ySf9faIGjG5ZExzD4AftVvaP77HSR7EPQIEk2iEE
6UYG44EbR9KtGPKXRUY4I0+OD97BYYdalemsUpj5gLBBUrWaN0cb4Xagfp54OZZw
cgQwupKANO42xSMRxtYd89l464MKg3/cDabyxTGAT7mlZB+ygoENzkr7hDFMge0e
XHkfZXAGFUjmp8gc6gitPF6AWILbBSxAtrEPBOH2YrGFBhC44cvkqTtjYkKJsOLx
mXTI4YSzd5JCEjtKqkW9tc0/qDSFZqYpXDjKbS98XOsqH75kO4aonvRf8jhYmCzx
aY+oIfe3s5b/W5Mh5S6hIm+fydnlQOE6HZzPbsE3UwH/nnQKjLQ7zwzwMK9KeplF
6jLIQTLUm91eyDSRScRO5z4tG+MoEXU7sanqX4KEYuo8a0cdaqrjFpCVYucNPz6C
8zfCk8vlsqitz7qzEW2BhAUqgGEMTwDLdLr0YcNZgLwxfabixIZMS2XlLV8eoRvp
HqGM146zVFib3yflsvoxXd9EiejcgAeKmqx2BtOxjtIl2YlfrpjKLJNS+2BIcSJZ
Qsi+YOXHgTC227J3nXBRu+CAdZI7lLcJA7FOxEryyFEzGvcaueS0Tahf66JCzSgt
nxC2gxRePWMgQBU/0WNVm798uqFOdAHofg8Ut78ZapWVaRNXifK7+E+rqcBh6T/n
3ccUcZq+rUNhtb45r/a3WjXVSvo/Wx41H/U+uPEii2rcEJM5Y/xVBtvCwUp/zd7H
zG1cyn36fI3CrpPktzsi527KlcN4NhzTJDCGtB+fcGWztE9qXIe414YBxyfENZuu
Yh0jz/620+DElahGfkF8hoWILhKsxq+B/haQAmjbb2ftTvVPMmBHYFvRHRtIlFRP
0LYleKDTdtZUCzwl9W/XQ6+b9Xv94+zR0UcmXC4pjzdPJeZ5rnuHDaOvS9dkYK+C
52Dob89s1EhvCNRP9NCN4+2uQvIWhiD3p9G6wlnF7+oQuMJlQDX4oONFetlCjPQe
leXaa5mI1/XrI27Bh2Ft7dpeC3xQ74w2rrkt46+4YOvCpbzzEMf8qzA/fCR5KKBu
KcMCvLzRrQI67F6/GjvUevJxaJZtbicEITeggRR2+tcSwh6s6hH/+P2+8MG++LLc
xh6zERP9BdBtDzg8zIJ8NjyQMtXrcwlERwy07HwtbBDfpNHecncsP5O2AKLhqkr4
usXMwvWfGMkqtXwtPf+c6VbfgPdD/qjBsZ+q84Q07E8D0srno+fqrScfVlN7yDKL
DEVWN7t04f2dYPfMZfuTvZDqHsP5hPnc3AnybZ99tf/G6rmljjFDcJZnK2JoD11L
KbWn/vUDZPGxWsHQYNr1BSAeZXzeMQgcJ/WiuUPUS495RY+04psq8cak7JHvsQB3
/+cVAg38TCysPAIwG7pkjxnwLBPG/CJ6LWYYCVrr7VYURIPOrJajbkILPJgYB28p
YfkFLpZYMJsD2aQ7c8JbXdudfDC7gpWDsO9zeHlv7kCwBoQ6/6o03WDS8zhEYJ9d
RPaomKU44AXxt/0JQHSxZPYH7m4LYQsxQznwgaUqHj9YzfU70hRs+zS15BRPsaBe
hPIsb2il3SEa6ItmBvWz6gqA9SRb08DEXhtVBEwAiDv2nPE0zEfmHGNzXX21PHWd
70P9sM3f2UUBfSrVNKnsh8MVGYYrfhkyUoJoUo2TvHYGBINSWgMOZhDnS1JNfKrl
hToAvDVktZYz3q/GcXDb2B0KnstUA58sjsR/SwZMa4b0GQGiX0w/mQgMx8KEx15Y
Wma+9d5ImyZ8Z8QEfnQFXL7m/RGg5FETVKsXIrzexAPeomCwiugbpYXJhl5ZmMaN
QgYyibXPX/q2m8AI5jw8z4kkKTuZq7xnroMEFZakvz1MfOXAorgYcw4oc5NVzLef
wzNFutpgK7J/Wst8XgkPJCBe4QiaLi6r1D2xk6ftDMZQnqsrTuqPfg5MmHdGx1ZN
wyUoJvbSPPl8hOnxDYSN5vB99bOeOHKmUcOTlB1JsaR32lCVD4tJX/Y4rVwh+W5p
f+uNoKwmosBUQ8O2MOO3MYZEtXQJTfWl9bB2CjdQXj7AdPPqlRdBV/pyRbSeyAFQ
zoi1pAJRSvdAQl4r+C2f1XVqxOwMS9ZtVUVYiWJwKqDhEOdOrsS+ChYn5Wke2Fy0
oMTjMv4CQR358YuUjx84b1UWCmG9q9vSN1bIeG25K3m8XhvZoMS/SiCjFb5ELye8
8Shynu54I5drpjBPbMIArHrKGgA1hE+BzQTQ2RJm8lTmhTzwqwaDgqTkReY8ZPPy
x+VZLjZizWUyqXl7bnI1EucOjQRbd/r7sTDoHEjE4QJhD1c/MgkrN0dwtzBNYnZH
2IMSbbc/fz3VU6nIEixvfHA6da94y8n7tNMg28jEFTf677MM08psH5VPdlhaUVNv
xJMCCCXm2qj3KCeyyObBxQUb4FI8XgT89UtOqGynStB4/Td2Rtc8WUgxUZH4SV+9
19bWcaWKr9wcSy/aOi/8dPiybuoT4Kn7ZtSIC8pkpSd+qIBErAAt/DtC8VW5mEZM
mVFE/F9mC7F8iITta5CPO6w0uyVgA7zy6q1VWOIoPAdQWjh4QR97wjVdo41uozKj
WPLLQ0PjwRRmtAdpNaHK/ijkwYokXYq/y+dXPQouJdK4mm1cpq1oVUxcHXdRrcvk
QK5YzD7p+y0+bD/+HqJeH6fxJ+ZV1MMYPP7dqSC81XAEQ6nKfILJaXdTprDn/BS0
WhIOU8cAqJ+0pkG+ZQhmt6UHyME/eTcvbdfAYNwaXVvk5FukN27+Wj4jUTCfJqxD
rGCl2LXjOqeVcDfrAyDWFYG4CgXUKwbqwZAY6aVqCRP4+HuBb9MELvJBfmmbEDO2
2YTjFtJa0h5G8lY5sB5wAgFynI5qpp+XYTJEEIoAxIjWvoAOhNwtTKTOy8xwGD8D
olOjQEmylBu6+OwWY2I5DB0CEV/m/0sh/4UJLhzuYUxGY/aumBiVhn8Wb0UHya1D
wB0X5qlpaaSGC7cdPO6juyjzbwqsgpq+IbgZ59lOlo4T99GSCPJ0laAzLb6Gdi2y
Hr9ME5md211QxEVgGMzgZFcea7BR0abKupF+nmU1NAbcd7BdhEBBHk2BxuWb5YFg
VI2pcllZ1+CaUU1thKI6i1vRMarLom5ahwFLde2RqWfS90x0+NVjqzsarDGIRzpj
og/YzP0cYZkkYeRXNrxsDngB1xPyW0gSYDTxiDpZW6pUjOfOYJbWvwHGjnOneZi4
ay0T+8WtWAT5AiO+i11JlpGN4UIFiPrEsAfFON8G473pyG+syPdL/aUi7lrb+sD4
njek/tLa5zUE5NsKC4QT4o8bVyuH9Wr06kL+bHBQtliB7i+bd0vH8l/rx6IaJE49
OxPGp8/Nae4WpO8WEiHNJxGFmkDxJSQ0yMk0bnFzbwVXdZqKsIKv49ZywDwK+ztq
1H3brY5fbn2KLSC1UwIfOSdbK/0T6t9DP3U65fvPUXPqdOdIc55fK0vJ2t9Qq5WA
DMmVuW35tSAyI1H8z9etFva/zGPeUV2kp6TgvbWKtrtiDpTbOCjr4eIDJw3IeRtq
hVfQ1qkx1eoWcEX76OlqHlxZ2ZqNo+t1iRmFSsypp3r7j6jyv4+PK7oDIQapvBgX
Hb6yJZD/r4Pl6anYWUzacF7/UkQS57TjoD76+D2nbK2UwzQitYFy6L9t8k8O0K9D
RXNlGf5Q0Zc/CktbsaIwxvldOjSTqegDW2qKK3/SD3q8Z7b4TCNU1n59NZnFCR6f
QN6J7XYpcLZoaJG54Y9EH4zq1Nthu6G0nWuBmxwYQUMXLT9d/wfSa6ymvDPt4yRG
9OYo2alEYHVTuNZFIH0du3icru9fOmMHFpb5ZVVdhLkBiq+4Re2vMdUT/vVXnQAZ
M+1i7poKBk+PCE1x4IU6V6MO1Daqmtq2wvUDGPp/o0hZXPMAr8Ri43DhdXkXjJpw
qe/YNQyigBSywgjbdzRFfjMGFzXjHDzIhEaL8L5n/B3NH4sDbZCTPGirECkqDbY4
3V8912Qh5HWocUqrVYdSwICSUAxmjS+L60GKe/9EDCXVqBehqlaU5pZh4Ddb1wcS
UVeOhRpqNpjLlWiVHtc0ynxUg/DWmHLQfo46oKZBnTOTEaF6wwA/0hKn2sibY0le
Apk9EZaxeiD/w6c54x5B8N/5gWTL+a6oPT0Vfv0yYXAKebZp0jYH0JFfieWD5Y4V
bQVPvYik5fU70WBVlmhLbn+4BplfnK4neFnlMooySbAX+hcT1vzOcND1oqStsWnc
uO2Mq06DQTB0cLgmQQhg3mRso8OBB/OIdUjms6RFH2uOcdg+FgYqpX9hgzN4e5zX
q4MLeZs7aJW0Hm0EMQfPkhKRPRntFAJuZ9zFJiwrPSDnfQ3dEqBkBRT3wUI/HMZS
0GjLzRaEJZJjFJlbs3sKMrAk60VVR3iZCYVB5Bla30J+8Jb4/KbNnQ0G0WwOP2A0
zeP7MPUhgfXbfd1mRMYIjrjScpJkWr5s3TSMe/TCJ9sr1mH/vMfYQ6dk72UEDIgw
xwJUJuH0zQ3PxcAwP4lrpGRO4v8LcmWxun9jAVSemRfglZlqO/DaaGTORxwxALou
yd8kIaI/mL8Axuh64CQ2jOfGrquO9eNncRK4vtepm7HZ02lB3A5KU6Wqs9/nmAYp
EAooDX574l9RclsctE63G6qM4N3gvXFXURX2OrRHGF2HuVH6HcgeBKktv6GpMoo4
M7OuI8yz+GVRcyxhDJiiYX19PLwstDATMZ19U173mjR7fAjW14e5L5LJwK6BIxDR
9C/X62mgpcMR2it3+r9B45NQNzGB6Z4Q6o5bzlwsqSjSyQOS8tldMvVcGHFNs33M
ltJfLdpd7zfoidHko1m4uXYZtqZKIFGVmqMP9rtp/a/CQutVn2tRSQw8x1ZfqTFH
hCyrab3nLH2y7mm94JgKTIPc/LmnKnm+H4jTfT9kYnxITJoq0r+WxAH2yVHN/r4E
T/uobEXUT04Tf//FBzRImuk1axINJ5ZWxVoiX16mUfrXoA9bNLugzZnGpPFm+LLY
QIeKsM8u6OebN81S+UNE9MgtmbAjfLxdI5HLEcEfCYbEArmJY0YO2GzWCV1pD4N5
22qdIMldo6PUzt2yb4wpHA1F/fKRtrTvn1Lb43mVp0xDD1bMoBAR7+h6PBNTX9HX
LiFiG/MkTyjjHlY3pt8jDTSjKlGYdfZsqgwXS7WQ/Gn+wh/gYoOsOan00Jc+T8Am
rD7M2WR/8t+We0R/vIIykgTvMenR/J06Ji4FD7nDODm+/5l7/Z2mkR4Q/HKRIa/a
dsOa0vr1mdTJkEmb6IqVO5iL4CYvG3wbKza+HrMAO9rowNKE4xXUB9sARStsjv3L
SxVhMRpDB1fQEb9e+n2AmN/6W2Kp7yGvRTqL7eUZXSZrl+aeZsEjfbYGhJcL6A4d
POa052pUiKOg2I60z/5GO0rOU+P5ixPlxS+jwlgCXT9H9gPrbbD4xxwkx+iTMjzp
kCILX3gBe6/LrxKoA/ebvRmnXIhkB5+PPMfz7J81HrC1qk0gEbNl4oPAcqtDlz/w
1R5AeVKK6DTabyDE2g/4f3veJK5qojIIb5+9DJSW2UNWiqxb4SITzgNKQ7KwDVBY
gwQGbYvueYk3pxgWCVvDFbcaRn8argyZqk3ZYUqXZa6DTzdrSdKYMTQZp/HP8OX8
6EClWCv8DZSPJ4t6Oq7AYCYQ30wlqoJ//ixFx7898tW1z5KyyB5q+Y66gS5ZVf9p
plojBcxyD+jf7YPvRn+r1SMaakjyvl0rE4rp/P92UOEhS4JDN8hjz84nd8uqIG9a
beI5ec9121pbwFWUL2Yytbn+blgwCQtvNyZkQIb53e2k2hxJG1+qvBy9TuZ4suLA
JX6Y/aQiY1XKM3D6CkIx1Y7OaDSB5LSJVVieit4KIiKMjRx25UNTOAJK0B27n0i8
YpC9pavCsPjiQ+xygJ3JFuTDWYY/5PHvWQBudOUpYmHEom8emf2XDjeUJXs0CZCt
mPerkKRD1zgyj6mevOPjPZvDqh2enYAr6Uf4vmYUypHYczOpUGfpcrIx2ls1wWTG
xzYcoA3Vtg5efEyq0lzmCe0tSoIBbnKl+tQQUZm0E6rugYU0UOUQb18sVvvVBtWr
dysYcfJDi018ECZSoe4a7U3ahSn/aVVYSJ+0jLLRP1WxeLY2oMBI7S6Uwwge5kRp
m673zawHohvTTX4kbELjRhQ7QIKnyQqy34jxl7l/8ZEm/9CvtQmjdiD40RU5PoLJ
af7dGBvTLI1PJBEG0kzmdavUoGKs162wEHpgD+Y/rZ4NlVNjiTXUTj0WFW+J2Hbk
YFMtPmSGGZYU991lQIB3RkSggOOfVI+iaKiUkK4xhZQEyM/4IPGIba8LViu/Y0yQ
yomFGbWg7FVvMYCrcZp1NWZJlSNK5Dv0kce8O2BmkIP1w8iwXYGqzWdD7sDFI8wv
KV+kg4jHAmjR7v7MS1q759cNTVoA0Oq4Gz6K9TO4ouG1LiQ5e4E6FNXSPIIS2mrJ
gaRqpoLmjYLnfiXz16RG4259LbuYnDFqe3nrEYuAB1h7c/i4TmuJscAAZAoWS4Rw
DZfNOrjOZZ8vI/MBckrhjxYcABnD0yQEcfeWTbqIehQJOgKc2a9tcV4UMu/Rg+Kg
e7BF4BAU39vDHQnup9tgoa2Txlo6APLLTWqmFGsnkNlV+B7RduCjMlg0ntd163m0
mcUtFv19KN0pTE/MvO5TEKMHVTo7ngVb+ExmekpfCs4sWBNdbDFP3+DdTSn2Avqz
l6VAanQNFXcafDdz4hb6qyKriPaIsPTz2cU/FAd3rHe9ZTJBNTOC/TqD2rzgveJJ
ULAThVo+hPK7pGf67hw/r8F0Ek+C+UpuQKWqzRQq1IGXMia1lw7KHz7CR4pT/ZpU
LD+ZwXgheLAvMgJPd7DoeXQNm+wRB4THskBf9yx7r8/EPjP8xClSpCm9DtvHxznY
Hbpf6OpeSkBu/drNSIgt3eVS9k4l5rn+VqmaOAqhJt+lc0EQTaR82nIlS4CE/Lnp
6n2M/3TeA8gtfjqrif4K0TrAU5qTk3m3YzyW8pbaF4294VTh4k4LU7vH7FaJYdWD
trawxqfQQz2C/WAaZSMmUejmF+FvVE7ArOOSmSLM8wcQpjWrrJe/mq77kPKq1BxN
AzO+cCJEmy2VGHCoXI9gyq3pkrCt8a7x6ZCRsOqze5vR6hdDfsMuZQX2FrGkFGhx
WJG5kYkdLcLjBcPmmh9a2LaH0gIvNh6jTAOcm9ABCzRmo4PuIzRD8o8kiMd0z6+/
toSw+AcszDqL0ELLi8Srw7mIpghWnWMr4YoPYb15mbMrNt43i1dmvcXPGvAvHEfO
+jrQ2PzcP7bkHg8ZL52zXDgg+svgPDy+6Tr8mM05tD4L5PmJT9I8XfRpZ8M7Jw8l
ONVbmtaShMHJkOUxlABZImHOpCGyVECbzxk+Qf2CZ6RLNpfy66aliYMJ8FUjHQio
ArdbAoLo/O0lfQS5QXV1QMvA4pOpBK/FTCzLzgFkTeZZX6KJM1KFkFQ9FeAIj8k4
SEWFwz5vEl3+9DeQcotHo5LJ1UI4ONoIe9/uOmZ0mU8oZ5iIFRpsczMZc+TlDvMr
U36DjKLgI1bsWRROpCg1jD43IS5Cia3kMwj2Q5mvxh5FIBptRKwk0rGHVI4BKgqW
ftS88o22mRJ6iymq7pPOyYIDBd7b2+CVicP7EV//BXZpLaca5fAsiOyhIgG1c2Cv
UtP8vsihwbCGBgTggWu9ZKlAXJ1O99x70rSuXirBZ38wNpgpkwJDq0Qg+bPA20R+
aoXmFTtB+RagNl0XIU3H6ylI+S4Epo4llMTQ6moBVUW+uNLY2oWvL0hmoXAqageG
Wrt3hL8Acul105tF2Vvb7NGtTqAdDOO/vIdAGR/MFDzAxtDytxfdY9jMAMgbfG5K
DVBLfsBqKWi2iLz02pchFB1yXPf/b7u7vOfbd40FWJ049eskdve8b+lLwL50KvQR
yRrbJpAhJ6DlKb9paz63BjVZWlC7aQIu3AkmGY/rnwuHZQReCsJkE/4RJzX0mFG9
MAqK6XC1i3HHgLbSMHcv7178cOLgR5ac0hYH2SPKwC25aZt0CESohYiYMqO/akWC
+CLOOwtKc/BZP+kD5tkAD9pgSF+19hoAtPn6Or2ihA4UP3Zuw3r9z4rsbkjXCGnD
fLc2IBQUywxUQKHikr2YN9/mrVgGyJ9/n8SKFIwFqs+aPmgfJDiWJ3XVowmQeMzY
3MhB/lCJmFZrJOcZZrLZuVnAixGFkcc7S27tTHcQIUN2okHvZJ6yrSI24ybdxo1f
8kM4Yk0gIAr0Fk36gP8fHIoH0/V19wlhiT1h1lMAswyeg9WqrVFfS/wF1i9Z++Cx
BopckaVlPzls/B9KovSkxMophgNSodNrpBXMA43ZwqtHX7UKWNw20sCbVw2m61LE
hQH3SFRlvjc7W0Z+G1aqrpMfa7dkcYZEFfzZjWQRK5vIm/kwu/OGLXZfp6A4bPoJ
2XZZRxHmHEKV1E1866R8kIphNA0xw3Va1i5tKzKhZU2SwBChY14o6V3lzfCmxEr1
MzA+bSLl3GtgPhFL/wpv8uq8VGhVZ/D7csfMI56TOyeCWbIAx9uEc4ia0Xhq/0Jw
wzmqq13eO7Z69IEy4lmOQCrp/K0u/WO9VNcRGcreHRDhvTxFLY0na4FZEY9EdZ2P
fAL/4go/2jB10l2JCEZNuTrGhaIPuNOg/Cb7MVwtWQ+UuCs3L2N0BSbeK07aNSnB
+5ogYbtjjiw5frqNAnleihz4IA1juaFv6AARL5pDbpZoRVGK379XszmoiGLK20KQ
Nw7lVqVUCN/i0N4vjhhk43RcylQPAlUnde6icp7UgRWMQ2MguDGbK/dbTuTOemhv
VjrhauikLyQWhCq8aD8OZPVkgidUSu0s1PKUTYcT7talBM3T4OFBw+MoBFmIuism
ndhdJgV4VnvRwm7L66BG0kGEj0qm3+Q/RYZCVMd6FeZY9++rTWkrCrqZQDS3ITgq
a7Z+gtLcS5erL88KTq6UnI0PrddTBiD0PWyVUMfcPG+zKgoudI5CSuiQeiZe/uNm
Pqmwbiv05KnUd+M7r2npiIWAhCeZ++DuIeRCnF/5De7EaEP24zYCoEpdjHHLUKCk
1z/miMwhAgDJboCtmFIF5sBMg9zJXYkU/JWC6wj4Wh8ofgIFq4pRYTvPQfUncAn6
e93XnonTle2suT8xi1nITY+2OB/+BsJbaCjuK0PDivQLI4wyGFWJLCDpTclFhFcY
a78dUBx5BD62DEsghEH6mokTobNTNsBU9CSQkOcdzfEfOpX0Gj1OJonYbqk2WGpk
mhjAlJtXSeFNIUNthitTk94TfxkU2D8SFaKQJO1N311DpVX8zBGHBiP9CcastuP+
kn3JJ4NEl/rKeYF0TEMj4K7spcDpGPR0olzxiSKsRXZCR9lLHgGWD6cRm8nc2t7X
FZpUMG94KoEAem7E+PtWI4EVhlJ3dq1d377Tx1+FO2HjdbXLpr01JNpsFTpy/TVL
FWjIwJ0tmMEvRTME+yKblKCzP8s7GthMJzogQFz2n0uFEmGXEBerZLKmltnBsP7S
zyGpacwg+XayoW63DFzSRk58IQwR8ohLTjuvM57WA2wO2TH+xiGhmMxirgqpH/sY
0Dw4bmdXoG2nzewzM4zhucidxUru8JLE3DIASCPbWTqPnma6WEaLk2QEmeijgu7b
+C4/s22gRSYbMtx1Ng2Bx28xywZSIrQZq2Gf1Ogpvhfz0bNStsySBZ7PA87d19Bg
9TK0KtzPsjeT+rwB1ePyjx5R4UEH8g/NLDAI8xYMUrzjsjuESgDxJEIrXRqVT8AV
MiQaJYj7hIQLICeKQ5iyyzyTUWagNgOsgXBf96cly+vLPRvg04nea2gCiiu1jXfQ
H+QCkBBdkbgvLweMTq0O8BWwX2gRLGm4EY2i9+Z9+SWYyt+212fGzklhxcgPu5Pl
J/pqVN9Lxz+HxMDUh22TecIKiojCLpionggMTLoP9RonzPkTDIRzGEcF28MOTmhy
/1R3HQg1Pbu7vZj+keboF2LqIv7d2c6VM3bEYywvdJMWSQ1wDrzYFK3onhr0oqQE
woFaHTIQ524yXDfJ1IZ3tOp4ql9jWYjpJWNdkLRIxVBVl5Q+ioB1ykXhOFNFvqst
FWIXT+UM+XXEqpKFEZ0SOhu0lAzBzXAXsriilkTPW1+ws3ZDSixWAOymR8ntH+np
dyWRNF0J6gRNaBl4bTBPryvI6sX1x3qL3jN1/ztuRJCQiTKtx26fKKU8KDZNqabY
DVO2aIEOMSeyYTaNnzEAjfqtNhc8mDW/GgHtpCftjDYMM0qKNtSPI5pc7qr7pgV2
a5sa8rMH3BDgnkdOvSQ77dk/4pvc8FUcylH61gGGRYTusg9I73AOd3u5PzNp0fXQ
m4I25UHDWjlEYOzEEJ/0mAN+KumweqtfkTlPnpfLw73bchMwtbsnjU1KUbArl+RI
E6Aksz9q8M3UPSOWad6ADnALYESzIKZhgNUGOodSbII1cNYwU3wDRIPp2KomV5Tw
M7N3+YglUU35L3ZwB0ghdeT75sotDE8kyYnTUrYA6/n/I/qaCdA2u1CxgqSd/9sQ
FReIIiL0MN96pmnE0KGVnrX3bKH1t3ELt5yobB0OULC0FlYfINJ/6hSEoa9OgFUf
ov3njEoaKWSVDHOSDWXKRDnAOWQpi+CnVo1rlc6TSfiKwnEH39wNaLoQsSSpvPPC
qsVpiVYDR0VvW1w8Q9EbXE0EUBN2uIOeY8wT8thVAIsD3a3GHaHePHdo2e5kzs6O
v86hq90upGthRLnPJQMrbGUv/nojVuxDhHGIEFH4oFctzne0kHfQJ9rbYZQN9Nge
oF40W4HrUc7HrkBfESusnM4SUEXtirlPOyzNE9vtgt0SbNApJLEHWtfQp8XEyXQx
r2O4VnK6Q51VLx9GfBiUFF1JsUGMtPiUG3TosVPkSSaa5JC/ScnhAIKguQe9XddZ
4jJzAarsN1iBJQrgjKtPhV84ia2IQjoK+uQ1JDDPOssUL5diCjksgJZh3ftmj1CB
AkrPAzkeQ4fwqKky/OCRvYC/VOxEBIZsT5uurpWOLhdQr9YeVk6f5jBr2bwCF5yg
skNx8gq1C5RU5Q98drqEyza93ZksRJEWUxSRTQ6ao2gAvOFsyOuHhnNz5T51/bKW
IYXElGuVUXXjGs1fh9Nnva3GzwzaQcPonPWGhHzH/vYh5Wiy6NBZ+evh7j0JIpGq
trrJH2sAKycnpHHFt0efac7KS604AEhDIDQ80yLl1mYGCKxiY3sZy5rxS4BXMRhj
Z5Bg0PPdFg8qtTagUipX6RCsnZsP7bhqR9nrxaxEAXT/WNThJzRH85JVZg5gBAis
i/GO7A477T3We3xWTsiDa/2IKV+RvKzJBI1UmDep4hzlopRlVte4t7P2EXwOpTPX
iYYqIvEa1nF2DOXHcfw7bL6QDEo44N1UujXeKf7MLfyZThNpjhf1RZYHV86ccSG8
MKJ30pi2Xk6t/5jEKnc/6XpyOM6/m6aH/QgS8gnknPNDWHyfwSyJrrnt8km4iJj3
kHLASfoAtSvK5wCLscTagimaDaRRZ6uTPMPbvWl5kEp1qmMubkg8fB5qjf/9iX+P
db+fQML1DlJW/gV2cVrEyNCgjWKBdsDVYiYg2DXGtanNt1JQr/kjDrvAKiZsApD7
p2AKERoG7cCzK+gbP04YxNvNcRfFHQTIiezC3AOl5UH1vxyxzpO7/Z5nb17RXOKh
rDQztbm0GctJw4mUuL3KYdjKdKroOt5QPMTX0XZDBZh0/cKglsfclIWnwJ1mHcvA
Uh243HJHsimSsd3T8kn/YD81rRDfikOL/3No5O1uPpl9zJ471S2PviEkSC44rMhE
SZOE7PWBBortpURbvtws09Ue350xqBvJ/VKMNwFfzPWKMKRdhxDq7nLzVKb1oBC0
C9IrjLzrM+jD2WK1BSRSEPEn2YHWmdqPk8BKiL02+cBouFnD1R0h5Hb4u13mN1jf
zxPjdFJ1qjz8IGfAWbcCHyYyPNHy0A/SEX8G/Ih2rq/B/EKtcT1+kjihpye3kgBb
K87rZ77BrY+T7ziQlwJUBDr00UNrkxWhdVUkxPDlSriIgcRwqgjJ+ZTdEC7QIyE/
kqPLpZ6D7gK5FTChItHQSHMQhSXiWDdTAX/8T3myx0O2qRaMtqXYn+k0KM8Lo1Zs
66Eyayox3nr+gHiITG0BOJ59vFltW/Nbe3n1fvXAx8TSMGkuwRWimZ8drnk5jWuj
IE6fp9pQeEfWr7sw+CA3eXuuOynVg4+GGGcPK8upGTfDyKqVvUxvg4lRg0g8skjO
F47RYlC9smfl61tgKDAOznm+46Iz7mAFB3bV7nqkCbogdH5XzDVQoTFwB8cK3JEL
ksna01EeRxr6vhZuO4fEufqWQPviT8zSObzAumbrpUkC3Vbf349v7Jslxm0+Pt2Y
+lMZp3dbSjBb675G4AZYZnNArflvVYfHgLuOKowFNHS7z2v+6B0tm9G5Zkix+G2b
U9xoA0qR/C2fZ2qXuL2ZustW2tWME6gtABtd78u28pnvPXmHcwRuowAJhUQ7Ekg0
lrrNj2FEJ5Cp9d3biLuM6LumKzEH4pYf2dYSa4FmdacMrq/h+JFrvmIZh46XK2Ul
8oevRyOqx56hBvim5M6AefamkBXwxSPyJhUaKR+sKvM0ANmfeZNQku3JazVT0OVN
HWUTKworZZMJNZPKHtGgrsQKKc+4c0dhu2zvLN+Ub53OYKMle9UqYwAbX8i3oqi5
H3Sso6SdMJrkKWX+wPEITbm1aOw72tcSI3ohdnOGVD0T0xpdVIVKW3bEC3NDiw0C
CVRASzNioNvFCWylDGLzOGgC/Lf8aZDDmo+57onRDQahx7mB0LG0aNWzeX5YQilV
2OW8bMgklvRLyfylKJxNIo101KudzgSn8VPuzryFB6xtZhI5Hs36svtZty8pPgJg
ZH0K8EQkfjjDS7Fi9Ht1kb7lXCctO2J98DUXdExCpalGG53CObzI8mIK8mTmv6Qi
M2bQaA36LULVMGmSKX7Ce8j6xWBV05OxrlYZC3ohd1Ytb04+Jd1lYR8DnvDY/PII
DNv76d3Q3KdJDB71tD4KbNVwIchCNrP+zJcjsQrQOWlwSTFyLAvRhv4/w+0rMg+y
KDrvxl7lAvRZ450wjaoADaX2nIRblX+RDHKcGD/aTH+wj2PTAEmBmq5+tgXCZqpe
sv02+r/RsFBlqxOtWF9sm1fsRQ+Rg8r8V0NTDqjXaFElm/vE8Y+xoR6rd7huXolA
3HCOdI5o0iVSQvtgnevkjK5EFYFo8JQF+xedGBXlBLecfdsaheC0sYZcDepuGUZZ
vli34ZJR8DO9Mu9747W/0sHGkFoYg62hoYtQK4Tf5Nqb1B++XJCzmjBFaIVDhywQ
WqRwNc6drMAQOqI8a7cpEK4a0Yx4g+0+lBfmSlKSmRwPi5k4s9uiwNm4OKvh/t1y
xnIJb2GkL0sxYDV3ss9QZma3WrVRRCdQ5KLzWPaIoRhB4dxqKfoMoJulJhkWtyy/
BH60Ff5CwzmuVq3EYP1pKNhvr68YDU5qLTaPvYR6r7O6zBlVl8T3w90cY9avgCIr
d9UuxQcQE+4mynw95CdLZwBTD0i0nAaP/CFXwnSENyyny1ZRvXI+18Ff1QMVyjDL
4Isa5pwfFrAh1Ghjn2TvEoiLpreU73mZfH3jx8pd7dmJLpKE1MaAsvdKeRy66GPl
01kQ7n3PiTdb0N1avYkJpxZSC0OGFNtQvTP27OPrDLpOALg1nlA3zjYgX5tUeLKm
UUlVeXDzo4qe4w7WbkP4Y3FDho3e0VV0GU5ZLxwh1L1OOJfOkM1jmm9WEcM+dzh4
TRgL4gY1SmEeuRr1SDeaR68VoeM7pC4xuajZwfbHejfldCuukgOdgwlZz4/xxfGp
jZphLUZ6QZa5PDIZreR3ggbVPspCfKwHXQS95vVfnM6g7DUKr99kNs0bO2FvkMNm
ErZ/8lVvbNXBWRLzZhKmJ5/yrr7jplBE8FqXWf+mCUO+U88IkbhaJT2tXdiZiIoj
3GcO+RQcUQUkQGfxGjzOgqea6YEATuCNAnjwcV+GbfdEYVo0ovCyHz+lpvUvakQu
hjQYZCFNXsqeTVhJIM9susD8WsfpL+DfGel4ibj5FAxIevqtj52cyQDdxChPzVTX
G1ea/ROuBO/Gar4Y/yp2kDPEefWgcWABTdZh5esTgYtPedDrkgnMLnZREnPJOB/l
ueo/FuWK0vT4xMYXa7NZaCY4W/IBGgehmsom+5rAyn9WjNnTcfkQc5BUW1s1JJx3
zWUWpDRoVVr1ZzYIuahASdnqO3mU5a55ZQ6M4APPr1fGYyH/09tPz+li2FWDyLJY
NGBbzuLu05lbComLJTzmrX7/618BJ8cd5tI/IXcfzw1445DkmJSAQ2SpdzkurnRN
b7hJKyfqOfHWp5cgPnwwZTXmSfszPHY8tUa2n1jlv9u7NaMb+CDyLSzI4pmrm4le
EiD05Adkl6cE8sIplgBoV5qUpkn+0G4guKZ7iDG6xysEySuZAliqU7nrOGX5SbAl
bDYrgeRFnFeiy8dEmXLJ+DNhm9R/yK2RXaCihG1UO38U40o7t5kePyvqrmAZ7KH+
O55kUx2uYMgatjgMWyHWlU9K0m/i6H5v25Jd98GCKNcp1gH1iz81UZ1KWFAy77ZG
kBO3rFLUPSLntsyiLxxMoo0cxJWVXCOpqqfE2Peh0qymqEhg9UetioqQg2fiGVVX
KOqGrsQ5Vgxl5PByu9RdjauKMteuu1MSU2Dg5jVZrI3dextr1B7sPmwPAsJPwR3M
hoZofvSmG4r3Ppjd2SPW89jW9kAXEM0ezz0vFhFIR+31yRXwcpxj0X+5aUpFItIV
KwQBkjYyspCP8GAnJDOcNAbgtnrLNBM/fXla8WYsH0KJakc1Xk9DO13J8fuQdEYZ
JiKAtvmi+nTXqKn2QgV99VjSv44V+BNJpcksCWUrzD6krWu9/nFTQUVzwPrFtiq4
Ppj+4EpJt8HNaVhGZ9ZRguWpPICBZSCAcXh6roVSixUzzFEK2irRW6T9MuyvM41r
6M6AO8fgfks7CQVWonHcLFOE04deCc6EO6AOsKusHtmbAl8xgmgCsQB9fcjik5to
nJT0RTRS77iJB3tfXUdIsigONB9xBaDbOLPZ42UvLrM6t57kqiS6jlLACFJROxIp
W5U8v4BlkVW8azAvJJGJ5h9AV+1z53GYtdbVFI1VZmlFmtMdUq4l/+PqTcXcehs3
j1Ai29BnIYa+bBuwDZOqEwzzxKBk2RAYovpQsWI67q70PSd2YxPYWAxUi/+fH9fE
ITJVkAfgbXgf1WrT3sLlANxcHK19eDYJMREx1k/uloseI1tZgI33WgBpx74e+MS0
8QUKjX1NACk8LPi5QI7f1sR0G2F+kjgk3dmnUOzvaksmg3tI+7u+R1N2imKC/6Ah
aYSFBYK5ljzp0eApb2eSAKBh7YMsclMvReXPku/5XjwR5V4Llmwq7kqUU5p+CjDa
TJ0c0cnCVmCs9lPxeflCPkDZvrssemqW/sANP3bh/7+ZK+ZHoQ9WzOpRsrGDC+du
YS4nyK6GkE4ioRyBHlLrTXuXRzu+3zl3xntxVzqkWpZ7lYtCtl0z87pMkkS1WCLS
T7D5CrEc3Fu2vt2SgKpPi4VtauOdkNlwQOdoP4XQYoXAnbRxlGeuDqahw9oyGW6q
w2NAw3hhHX6lwTU4Rdf3m8hgwJ9xJ7UQTaVlb6dhMmmPjkHCzNupNat6urexsnAX
ndwIJK/GPFGkrMOcCeONUn2Z2cfG1iV4ptU9axB/J9KAo7qa/M/6Ti9e/Li6LSwW
AHGzxmj70dU8RCsCmmuEQAQw29CeO3tuUu0b7TpPe3Pnzg7IN9Z3E2W0xAUYbBaC
cs0oEe2nMKepe1Pc4yUmyOoUuI/w7QFbOy76esPUXdl/h5YqTwjtczVZrOpRqQGj
jsjV2b1JeXmsxIRnh0VIIG9VtuTsuumlG4rKnzc+eR+zZh+kAWwpQkIP+nrDsfsp
+g5jQeQQbZMkj8tU0mmqlZr5K6LbWMIRX39pvNLbjJT6u8VWe9cAtR2x6ILVSh4c
2pJ1H6znmpVstMnM0Y3tSAyh6PKxpMKoI8/jhCcecOBcAB9wqh81IVA79Asriwmo
C2E/3sUPtohrV9AadS5ohrTdbdDXcBIRpjIx5tv+TgWmjaZRoYVrzUVCZ51aH8Vg
XEx/XHZCPjc8Gao3fC9uNZW9ThmmAUlYKw2Be9ZUx+/jrTO8tuotsDGqoetsn1ve
/F8h5Uiu3LnEfwQ+tIrgM2JPqrFGzi9kPFmgh9NYtiXmgcS3BD3lHn6ivrT0eEaL
Yz+Iz09WowlHhjYh0yPfWbia2sJbhfJZisbU/u2qRyE+5Gri60RehJ2yG6AWiCZb
5tVRK1Eawt/NzIvmSoyMe2lKTftpL6QO6xLHVn2lhPiht1Q6smylYD1+wVm0G17A
kxdYP8ZXIcw5YZK4FMPvxCQb1EBnb9gcETerQ9ivRKc/hfkUfl4sviZrAIWZqvmp
Z44ZOJu0Dpe9xKxEHnztHBy0W2t9zipexwimqLCyVhx0TUgt7yC5sTYjv6U83ipZ
045alZ0XupQpSUrR6E+LvCqgSCbRVVEiSCIk2YwJz8l+JnNNVrGYaFbkw6cSXLdI
k3RL4168BFdQZ/PNcVvdmGe25YGdxntouinITg2oH5uqMMcpA2qVt0OZa1qRDyAJ
02P6c00eGqf65V6s0Ch8BYG9ehJCXBar4sdImnq4OM6swp91jmhLupqQoFvc9fsa
U8x9r7nlCzlPRDhqFi6WkxzJZJRaS+y3xdbWs4T4n6gcmI753Uqq7jb2Gp06d568
NtSQmTa4DwPHrrP5RfS1bn0ghw0joZaATBSM2LUnJ9Q7v4FYK42uuaxnH2CHNYlI
MoekwOKriBtCtFWO+qUX3Yt/IH6omWMrwtZ7c+9N3C05tspLr/DRIdY0fwvvC5Xd
hjc/ANocRQxsXtJoz8z75vF6ev3YAHB+KvF95b7MOcUrTToaiU0Rz9j7Ypl8Jsbc
ZGQlzRzYj4jZuwQqn9SuSYAecoCPLkL5gFxjEWxhhCOWoLHPsZ9pOvxVd/wor99J
0whEPYAsPZXPdaYhSGS7oHH5nQ6WJmXhCrYT1C5xADT6iG0ab/ddg6yztu6ecW67
PY3INk6vjaQJytW6FewsGqNmCpQxk5NLNNEjBcMyumZRdS45YtXQwr0+q8F9fLbI
NHNQYvuoCWI2s9d85209BtYnAe8+7kTw1ESOhkxR50iYCnMno1NraBEbvoDFylzY
M7PQZytVVgDETVeYsHisA/VleTeBmmJqD99OWvcia77CPdO870IACcO6PJnOrBaO
d9wwkhBKs0KN3CTi/kVwluwD8OfnxiUZXLaHi+HMH4lWlbsyhGpO95eDz5Eg6Em0
p+Z8D+BIiicDYF78+nF7aZEF/NUJEyXBJ7hj10XPAw+zpdc1lDYU71u7Vr6rbd2x
OpurdatAvytuux2BDc3uBKq4o3W4wM3wUPTuNMBGEJ55QRUEFP7f0qGwjiIsh2ZM
bstH5zss2RHcf3w4ioBBc84Rr1L+uqxjYv8Fuk7kx7bi/MUc2//V3QuzCzHKcidp
fzqbkyymUAEHVqvLRPcBL7GYb3hxmzT772FgrDT/k0t0LlXTHCHeltu1NFrSFSu1
44TznjAVlBlN5w0ysh9EYABBkywe1mBTplANSrfK8ZL7RDT9B6WxM7IvqPPz0GOg
F5Yvfrb2vJ2r1DUTpylh+8SbAzPfRyQG9rGRKLxmFn6oRtu8bJGb5004kuVht8cx
lCb1uJF+Qg5qNw7XOE2LlyZmkKFGlbJ+53cKw5yvaF93ptw2m41bjicDaubU01Z0
uu2ZFZYV/voJaYW3K7TpW2j51FiOP2xUqzzKJuZeDBcM36Q3xKNtMZRGNawxxc0L
YlbeU/sZDqqlP1LvCSoO/w6nTvMHkmaZewqI601n1rRp6Njt/zjU3mRP3+UNB05M
rR6w46IOKyo7rTKQVPZHV4BH8BR8Kfu8S5d7T8vT7OnKsSkFR3a360fKVSqHiL2v
c/TnkLswu+kX1lgukaLSG0NrPMiY8uVal8bvq8lAOt62yovvNr3nhma1x/mhbyOl
AY75ESGH7S6JPqxBcpqGgj6VF9W3nz1Z0HpZuFsZPBjHkSPt1Yjj6dseBTaT53WE
U+liCTRzoELzu6jnlMmbiHEur8HDDmscG/0v/7KHhz8g8KIVe1+BrN2X5BvOf/Zz
TEBuMZl0jBGPngNKLJ8+GaP39s/q/FHmpNWqfwWkXL0biRq0zERyhb6uN1YHH92F
NBo6ECGzz90DqaRBnVtU/v5J1KbbJm01U0jC+gQO4tmV+jc4atBu8OzULfXB8Hji
Gn6g9rdKIN74QrWGbLoKZ7MTGKmwFdWXc7KtKwSWYeH5E/hyw3P/DEFUh33aZ5U9
ret4kzTy0DvF93b+6OiELGXj5/qnqZH7J5WSCvl9wXTRSkaU3u7FKMs9+yPPethL
9jqPkPlJf9f2alw8Zm7nyxwybZf/SVpVZl1KbmMpc1LYiQJxH3uwFlZsk6d9vu2G
BS1H9ySqSjS6L+CkcoR0SA9bAsrCPDkuq+xFDyuiZyCz+bMJxV/EPiOEC7Rco02V
g1xfj0CRGwMx1qIV0Mluan1uLA1SPmTZ5A3JbckXTUGlxWZSwVFjlSyRSVmJCnfi
TIkOcNq7VmolIzOOdPxY2s9p+VwhhP/yAzoNbYM56Onj0lF6L8LpeeUmBKv8Ny7a
JA73gj30VSuj/M3sXuC4caMJqqL6S6PX48Siy3CKmUtOpbijS+OwvaNWMsZSPkZv
fkMVeGf1epHTgI/7/KnGIYkEusvtAQXHW/KSew69SD3tL8PDzEJdf6tpZikc9T3y
KoujOFJTJt57XD9tdTnCyipkM8tPdKg85XOvjWy8jztG55azjgokCmTeA5kYxUFj
mwq55NLbzXTTsYi585ErJ3XebV5q/meWf42gN5UZ/Crr0VoXQMkM7GglxbR72kEU
dUn1gwf+cXXxEHEy0ABgmO3DB6KNn107zB5KDQbId9NklYrWUYYM+E6g1E2IKJ7t
i8oBDJQIBm0u7mqefTEWa7f3UOEs0b5PYOCwhTp1yauIvjWrSPq2BBnype5FuK8A
hEhxAN2wpzPB45+2hsX3YFWpwuF3tMvkkO6qPC8eFPeqDcbFKn4cLZO+SRa4HGdZ
R5pA0qHlQJxRFw3Yox27eSpWXz+Kvx4DN68XO76tFzh6vGfDEmrp7uIDM0ACgIxk
XaX6j6BqhaM9uw1MF+nccIepxQDjuT1h+CUs1GcShYV4c7gBXh8ycb1YKE7p0Qis
xLDAVkAVLWiDbRiA+CAEGqo/bGk+wnOyQQnaXS18/7qZE5r/Ctlt1YAAFbM9F5g6
Ec2iWQSNjPsKnCjzy9eYd91h7wMK4/LzSXJRL2LWPrevtReL0ukZjkkeaJtosnAx
JaAJKuQkkv9StGcNeCChEyIajN39InYFcQb2S1jPxQ7HL1OsPbH1QEYWFdmXfM0j
yNCjozcPU549JrockaXvyZZZ/ENeJ36BqXE+YdAN8Wf8jY9o7WLA53BZAiOO7GYy
YXl/LdSfhpWaMocgRTdNk5t6YFV6B+R7xFlXjAdjq+Gt4bYwMcKsKmpekYqR2Xsd
CHu8Zy2OMFhgjmGfiXYA/4wiw/N0q6w+zfiu4fsDKR20dbIZA/wi0pQyrm7lNru8
mutbfO7ak8h+MFO7zoWIOTIwZZLvGYeKHE/HunqeWQ0jF19TlYb/SFXxoyaS/KTq
0nVUB9dGqo+Hp5aJqndbMy8RVK/ZAHqe8PGYaWqR5tVc1XgGut75JJ2EokpzXFLC
HfR9BcfOCHUmYpXUP3AZI93kjfnGSlHV9JoBPIvhicnmi6496UjDgllL4+vaRsF+
9Iu7vRaHOdcfcGBSu6PHMClZjl0Xf7q16s88IgHQo0zFfICv17+YW4pbVICJSj2E
dghERbQpiltPG0Ml3oGa0hwZbJPkZuItTRTKlx83rvVkLUno4USSBQSgy81FfGcl
+iXid6jgmalemvtRQfuU4X+niz+P6OrjIi1EmOWV8+NVupLWlNHt1fe3vsTSEYWC
PuWRkpLv3GDbt9E2pvkh4tYC1ta3MBuigEPBtuQ5BKBcgsfnJm6khxZFut38QRgU
zVa6XdbEtulFmEAQ/qxf7Dyc5W3bavFIsiRY9BTBOEFshNnTuX1NZm7fMRqxkU2h
xyX+/znjByaq4BDKGtsKUzyakaSneX5mZxmtyaV0AgFSVdZfNl/yG5Rvas9rbU6i
aYANTHC38N+SaOIJ+NE0hXRk5JvXsjSpo6BLUMGnrw+fBhZUqYLIFy8Qb+vUWzPJ
WdKPsTuyA1Or+XDt80jvjdbNtCHUYvVmPG2G1mJ8tYqiJIvWztyli5DWc4Uwm3bu
St8/3q9EdUgCVxJzQYlImJi1XMYYFNMxxYGnw5IgUyUO8OpApC+7MGQ72hBBp5he
fSanneua5x13I8wMGyBGuv6sq594TO9cxiKpxBEtyvbwlkvEwRcofFqVsTYFFtZu
zYrdZ7OPUmQ/CbG3DwvNZMAzHFrf1k+BRurvlVlstfnrBCsi96deq13HI4nWncbB
JH3Ae0nNRQR/U3yiJosJd/SDbArgVdHAtbOlSpKdX4pIsv+vO8pG9DV5npv/paKF
dsn/DbIKTmJoGgbdm7Y33GOT3OFkq/Q/DNYjFfvkHieS5A+BsVBb9SXpEQsVrp53
j2UhBZBT3iGn4fo/752+wdHJtkE4SIdx6uZqfgmQCjD+NjUAbAxJOgVahI4hb1Hb
SW3rySUpewJ1nJV2HYWXJmIJYO+3EqYdMzONA1uYyMFoAlXqHoSA6ltDbX+a10OZ
SVYy9quH2fUPgz1DyofORSihSkKdYeQu+TnOYjVm71WrVUKzr2t4lkbF4m+uKXXW
fTkIeRvucV1Wv4RPR7YQLw4uMwgWsusEg3DjxXXGNWGofVYnjuEcd6wPFP5JCM8+
5QjStq3TtjH416ai3KnjPmaRDH2PrPJixNWodmqqNYDueJqtr+Hlb5JXxicHcrK/
GJqmeDkuDvXMAXkB4tENN4fqYIguTXP0VzJH7GDoYDYitTEWs4UgX07Lsd4pAg6E
seA9LseZCnApJNmqfriKMkRkTevAHg3FEZZ7Nlerm6RuT9Hd815ZoHjH8uGy2EEB
tD78uDDIksVJlejS+9buwixvozShb5szVIQNBl4fme/xQzCDEKLVHTyJd/7sZbLD
gMJopXlonAarM/jCQ4y4hP/5Jt1ekzaVXidxJ6KgerY/hLGTKGTMTc65Df4/px5U
TWTSSkLATPs33u4VMWme/0vfhY9YB+STLBsiZcddOkP4NL5TBBQg0KPJ6f+ILUvk
VligWu1WK07HaNOVfc9I/5B1+kgy/5FMkp+HYlgzhAlgKmfUl55AYlQ8fnpS3g6y
XnexSqwQ/FIMprTOsU8lKpokdf/bCjJyvYjjx04LNPl/fi/4rO861jUtxuvl1xQP
w9k0ZYq8kjXWYQywiot8I2vVilBbGtt1DIEBppKO09iS1Va+d3ThZAeT5wMLK/mK
v699nx1RddLZGfl/SoIlanQc9h/8nHfoJI0YI78j4BqqeHI/+x5/BctXV0hRNMY2
zWOUQSyso9cB+1rm8JKKHfWyNRqfK6Ker8XCvXCBkwh7Uy/LsOLKF97eKFhbwuI5
qKD+wNpZR70FyS9S2KZ0G/hp21chLxLgoCw6byoVTzzjVjAObLknlJNzuLZt9j0e
QfzGil0VUUeruZCLxLa//roXCASpsKdYA8tHqURHkoOvb2L8OUlcJ0RmyOgRVBHD
D+lIydbisPwX2cTPn8fnFh31vl5zFUh5du5jKsU7GFcCmjQoCdXYk0HZzZ6vgwtf
qMQQGWL1Dv/Sh9+QGiXk2v1TXhLOmO1yIMRn76SnG4+VAJpaTaHfCIENiJ2AT/B4
nuf5ThXsMtitiO9QN7ul4fcrK+z6Bg9fl7vVgwX/g1MT9z/TzdnScoTJdAfNR5bc
J2tw6P5Igw9gy9xkwJFXPG8Q2prbJdBlaGDsWd8WhdHvC6j/MZTQyQ0mT3vfhS5k
G3yz+3i62zwd1RnQQo12IBloe5h6VNFIgOobftCt+fiZEXQxleubD5TJ6FAp9bXO
UGM6aQh92pvPCVmz5q9TbB1je+55ge3PJfmTUgKvXqSEIdtG2keqZmaaEKSJya37
VvXtmXz4v1GvFtZVI3fyfseuHaVOxVIfnD9xtFts1WAEVNIf/z4RpV2gqbLMajVQ
3C/eIdWW3p8yWLWCWgkUltmkQ3OQ9DqL3kLJqVjQ2A2oDUi3BFf4c7+6zZIWBZCz
atUAUPUbVOoYNJH5savNHNrEZXd+sICsDmH2IbCW+4pXNraQzQGDzjxssy6SQImN
rKn+10eEO4c2Pxbdr1WLldledpzAUPsZ+kAyVpeSOoDJ2WXJU5w7BrL+ZK0Bporm
/z8QTsnUVj9O1OGLvlpFtn1b/Kk8KENY6WvFapO+B6txIlThhLoLAnzIwXsFrlXw
nmDsD6sioWhp/oTmm3+AsvK70dhVUvfSiXQ+Lr1oRbqELMh5Q9Z1Cx63e0H6oMoR
/enqZHz887FFLgLAlNTFIm9c7juNy1TooELPsUPD3CoPrgc4XS2pAsZ+rEcOlOmt
jeeexh3aXe9UU7XXq6L9JKuhu4eVIpiRRzf8x4rCuXeVqorBxDft/Fn9V3Pg79Q2
cr6nENpmR4itJgGZAoc6seNek8sb8Gf/i3UBWGqXHd8HNXJxx2GQqzElYO9QGM/8
AT6I9UaQgyGOJdJNVZfTR+FONvMfIo8JAkwNXuUqGCuNV5eYG7bAvV+78hwRIUoe
Ai9C1aUet/OlhtbcfIyAMikOp/Eg0fyJYt5niavlGYQImnbgZFgIdRzpPZ3ixmhO
P8umNJuqIHGc6hPD+q2+H4E6Tfpg1Wd6K6TSjO39khI4yT0AjPbHEqPthtrKR4ij
RNBVPqpjwT8kwTKRIZQtRxgmn6bew0/3XGc4otVpGHnm9E7G7ensHFxgAmyuBlvB
hQCqGpXR+P0AX4f1prduDgM5DzL1iLThEFaYypYJxdPfH1drL6LKAHNM+9Xhbexf
UKLLuHLQ2FlmfaF7Z7+AMDVJsePFxLLEO5R5+9tgWw7IUcR3DHjMYh7lzUrHJCuL
LhKRxGMTdsoxHQ2slJmRQ1RKgVCw3ZvfqOwpXdDRyh/eoR61/fUaGWFBuvOUGDg5
WOpMSUJnFSQEXfgh/OAzc4innQP72uhTMjcY/zx3UNDfruJv98nLIcPPfiHxXfZ9
Vtmyqx5KNgIf+LjPN5pVEEHI++XC3kn05XzscKElQ/iw4/cRWkNHzlz0QisZBN/W
LMdlr3qmhmM/zJYj9l9CxQg30FexWALEcNJ4Aqzx1W3bKr2MI6QfljKIUqKxvMYO
Wl1azrmjdSy59hZleeusm7DdwB+Awlacljkf5fFjTJXMyjil8lBqdduae8q1b+eD
jaWI/9wd50I+V7aKCiKTO9mT41gpbxHaJGQZsvHzYu9s77dOlzIV3kbMTOo4ec7E
Vh5ZSZBHYQ2qOJXqyTGwroTzsEtce+8UjkItGz1iX6MjjduKl8Q4Hwu+0KCB2LdM
2GbhCNnCnADrj3uo92G/b2iqz6Tuf03+xByjt5i9AyyQPDlkysJSKLHFL5PGIkPI
PoEasfylaZX5D/sUC/ju2adVGFQ2dtcAuZBiyBSWJIq4BL3syJ/WuigLUJuhGxRY
vUT8BSWjNkPuWoK2ZLwmYAjDFkfv0O+/WxVznsL2RbvgBU8nOQERKJXvmakqrf0U
SfAhZc8pLbnq8dkWzYNv5JNr7pKcD8zHNwVU6kjTu/x2yjv56U6P5VzCMuBE35Uo
49wym+bCfUxPyUkdC1y5OsG3GDepoK4O6t1sxNT5fnNZ4KkoarE42sin3YdCsII8
4Sqpydjg/q/qicxBRYn60aLvsYzFCQLVpxRc/6hsmJHQKF+RJQOgqhXfB0VBUC+U
oxf5Uvg4ursbbOdltB+Xs6AOTpGoBoBCdqgWBnl8CPjqN0q+tzG59HI+kGWBrWX/
dMe9XDNMExMJqV313+N7yPEaRCDMHM1obyGMxY3Fo2BSTveh1dwSl/m4pgethLyF
lEBmw/kO8PTKSgDddQpXIxRUjdT+P8hL+63+nNtiDiGHprmj/EJLSxKJqDdhBUl0
2UXwUpbqwkrk5eJRy2qjdhtcU/dcaQAqURFZXDZrW+FXLtaLRE8uYm9vgASnMJO0
X5gmKEBA4ZwIcRxqlCUluF1YtGMRMbbdnJkpUmqJbKmPWHQ63CGumnqbSOKI6Gkn
il/1CLAPOnw4awgTpAirh3lHXXUHJjhVgZp5Sv5jGF3SWHmUlKfogx15wySPkNzY
+35M/lfZ9ITPZdHfY6IbOohWFw7+eaKLTH1nLV+J/iQK1MHKf6IfIoANAbtIN+05
P434pH5F86WjLJUeeSAx3+bGUFSLFD++QfpELUAwMAX36gMvsk2WvaEmTexMv78k
ecoY01CZvJLbtwMqAmr2fejvotIkKo+51bkzB5X0wVHmLLu3ivQknwBO0cVV2wz3
+RCrbHv2Fy6Of1u6JTcSpjcNlcfTQbdWXNxHIKipgEH5EA2sCU8qceeqbCGVl/OH
6A9SD0XTkLU/sZ+aXV+XLrnEoThJzuAtM4gxnr5Oc8HOgLS6FSlKFvCgNIl4OFQ4
WKioley1+mhlZRDedOA1qypnqACuxqSpJrnV7sqrUOBQM7geLBu3tYVhF26q6a8h
67LYbWsg/ay54ZdrlazpgSGoSsuJtOcvj823hvRMtCRAXWA6Oa1kanYFGzDY1Mha
D7vKaQZmhiSmQ5ZMfYViJmn+SVB0l0H1SXo0xbni86w2hRwPf3qny7KVwPGcsYMs
hnvvRv+NievludujwyLMSev325/O4rgjfyOGSE+dd6gKpqZKNIib7/uazsofCE+r
iqoV1dS5zgRuvigpPG2UI292/eilQXC72CIZLBCi/xi7MEdc2ILNxbONSJlQediP
NVxL3UpvfFme9qpZun5Q/dwl16MfsljUO4/mxC0hvdjsjMnvgcTk3KEuUTAoN55w
uXl0vMiK+7wsqC7TUPp0QCEb1OlkoC6oP27ReTDpgZUDvrclqf5IEIQhKGKT51yt
9HNnyWKLukgZHD+Y91N3QWV0CF4LM5ZnGjTauv7+wdQedQbt1fGFeG4+0271XSzW
/eR2yJnfWTT2EvEl5jJyxhCALK3kXedUbiJNyY/qoNQi+rhjTm7BpDI05SeyJbfL
oHQw+5xdllnKidQM4+8m6CW2hBGhWde54DZFJWCJRFu0vElnxQt3qSb5MWWNS9+v
+iDcoh18zwjiBezgdYcGcXXhu8NPHZj9mewy/OKlJDu02OkC6jvgMEORFXDdn9oE
exa77S+xNiDNK0KtbE3udAUDVZtmYrme0RatsFt5BCwDbyWC3LGr0yVO3w1wnKru
Mn3WHgcPu49xE0UqUDDyQiRfsHD+i/3Fy0A9ssQCeUAxqLIIMwPJZE6xD+keFbyR
aw0wxwDbS5dBLonq6hGSx5OZO3Q2nH3MkkZBiqNUPHbkFOkl11oyIrLiCUupFPBG
MjNZoaj+DFE4vsGWCVKMc4Dp0spmbjv4wtSMzW99xfU9PEXDF8hugK8GwvY6dML3
bnlN40n+0MHkOW3sdovVg8UVB/ziZoxs7GgMrMJiygV9EOYBBJ+Rx1KuPhWSoIav
aBeSzmDpQGg4mTdlFCWM7eolaenIMte1GiaxE+c8KmxOu9aQwsx6FmSdBqASqf7F
4B5DfGfgqsPpPXlBa+GO4ypytK9fMxYH9B1Bc40u8pHa6N4skp1NfXmcG8SjrEOU
fU7PxKu5qGasS5naxdpL5QfdANtOYvJirufEt6zaxJFhGZlvzPEC/OZy7yegN+WJ
fBfUQ0Zaby5YK/XRzNaLrWrr+JrffmoDQN9jSlQcZNHMIj/w3YC5e6WVLS9Xhiaq
0865Vx3EkZQMpHe7bV63sRPNkXxksD7ggfo5hvjR+PPEC7SXPtOOG7Vksrqwrg/N
ej4R76HCdBsj+BZd9aTHmWv9o6umIqwbcPuQ2NsTAehKRz8KfoGT3grqwm77QMQ4
A7GhOFE9n/o3ADnImNeBQYgz/fIRILBIi1XSShYUNIjQJCxLBFrq1iLOA28GPLwj
yGDo+av1v7IbeYZ1osyJUCtz3qdowCE+4kXpnZ7vv3opUHmnjo9ODv/MhsNGH8k0
yIvILQFVdjofDvWD1797Upi/XBqEIi1Xu7sHEsMK7L+iPHm9Io6Oly7bYj192FYz
j0RvuIFxbxNn6DAfA17KAZmgopQwfdJKG6Vts4MTY+MH1VyOA9vkYPqEGPbr3/Lp
0cWF/r6CFQO23Yo/NIwKQriNSWXZtdNdFNr2tLyxPblVwdIK8KW91pyMZ+ZGHxTP
IUvecgPhgOsgKhra5jGX+dV1nGlpu4nRdpwiKWCBOBtBYkSPf8tvyKtD9wkRXm+N
OEYmoe9JfbVWcomsBEU1R9kNh7TO9ekZnZxnes5YNMB5u5Vfqi5BiipeLI1yZnmb
5qIrmxqos7AOWtVlIJosadzSO/NFfTfYXWx4g6T2bE6spBp/g/2domaUImW8l1L3
z63bvL2C5jdp7VekXWuxJIdRU1xu4ieS07s8hL9q/s6LF1Wo//4C2ioQpQibzHXy
6X8U4OukdI6Za/L4xODK7KnRpUNVFO6zuVgekIC48P6bA+Mx/qBMx6YRJTsBy9qL
qsa4tNJ+YNoCUjQ3K0w2n/b7Y+CLwdZc8x7h25IkYP7CTqTjRP47U/+UlGGD/bPy
ChOljsOpEIgeT3TZcRyQRVv8nQfA1iD/VOfdI/0dP8ljysxe7X8+yc5jocepnBMu
jgB0I3J2LVPNsnJtKN/rn1pi0klgsnBvTQBUOgH4TL/KVt6vT4A0IL8ivOYed8ac
3KlMLyZ1yNHhnDMbNDSIooRZacXqMX164Ts9ia2uOPDPiu93XAqxG3PnDy5w+Cct
RSyPU4LHXCeg3PXTQcwKML6vRbgUyzeW0RXtRmQ5shmrlixp4gDJcKHQUK1pQ5ur
hd8n1S1OVOqp2fgPbSIpKd6e+2PXSWz5Wcgy/pfxJOry9mvUWoYa+DZdP/irAHjT
xEsZbpadd2fDIZDFrWd2V8HMig6TaJhk51e7bU7Mf40NUJSMsYQwri8gGEnDi/zy
lYAucSP5LRiI9psL0Q/6uEiYCXFdsskCmdK/2+v8shupg6HHZ+oK11oY2mmE270m
muHPiLMU6LkRIgPt+rIjMIcsbZQW3y83VjFbMrHyPYF9XhSeqtKcqJQzBc+XVXlw
rVbXTTUQv5g1mrqN0TQ/wuZ9aR2E13ppbKcFAqKipoUlCPl70NA7gWDbhpzY1XpO
E4G0yBe6NRiMHvI70VWD9o4O0OkOPLAi2rQy8Mivr1/RPDHv+sXgX7tVX6A7Qq0Y
1i83jh7/eo/qbz3FwuqVRpYWbknRpP+KU7RAJBdQ2gkBrSFI00SR6NCN9jcdFQqn
c2fSM8ajw76zmjiV2qxhgf4ORehSHv+fpQcZU584+jAxhjZBdIbxnNW2e+VE5IU1
e1dsxELyjkAbIkvcKlO88fgGOBlRwts2vgYh9lkLEe9Wsink3oQl3K/TxVR8oke0
w0RkSYHWZM2ESBZhJ2r7ezFaxHq0t3DFC97aLmz0opeO3vBZh32odfsKGIo/KZkz
g9Mxj2+Z2WUh+4ObHVtWbafoqzwD8Qov4K7GjxLHNsE4wdkzZulXcwHksht6R3H4
q9xe7VweQjekiOJm4rwfuCjDlvih2KIi2vHIJsROVpJ9TAQIJ2NAVZJgWTousfgm
nY/0i0lH/q9GiQmt43k5IJygnd3d7Nooi2Li2ZYw+K1GdpKyrlazIGH9u3qVA9XO
87KIWN8mnKRBa+KwpCYJ4KiQCDIHchwmuRra0ttwEA9ZpMJvJNkClUdt8CYQoBDo
WC6jOa/sKkAOuuR9GJkK9GbcQAyzSq0WNQEtqdA1uYEnTmNeYRl3zOkZdymuGnns
RPXvimmAq2iqSN2PrTqzXx2ogOqAYJS+1bIGUVQSDJ9UmwlX92b+HeB0h2UgRZ+b
MDlw+DWhJjaXvU5AMyIgNBDpYQYdIloredORCWDSSHbbr2bxmSVHUBOwa2o/q/nd
H05K7CQ/jLlFOvkTRiJXMS+rP6FoO3DFSQV2XDg1hBHvBtRO146Q6E38kXPbt/X5
p4wn/DiW+5pEUM0DqrJ7dD3CAyNVMxEd7LQSg4qotdyCnyoLd0KdC+V3+HCTv4qQ
IxvaWttt5Lkt2ZmvnjW8+Q3o8kWYeORMkIl4+2jE5RzrQzjM0vosQJHtcuyCrFqw
LfMidHQayJuH9HPCnH0/MrISeydvLUmTL7t3wa70zcRLyD9RMrPzGqqZlbMzVtBd
r6GrfWtMEYaIqrBhC3JM6oMYKqtNAAKlGwFY4NyRJlzM2s26NaDz0cYzOWZxuGyL
qy5GzWPZpFCG0GfmEC4MBpO9cd2wA6tkzQq68NlYFzuO3DM9y3sK0SiIPREVfXo9
04eUWe93mi5Jnmfbij7+uDLjgJ32m/1HmvvW9j8iT5mRNUhIyj71lwbV0X1/1UcA
rqkPfibaKXuSkyKP48OMMWEzqTcTdSujDTROJ7A8pKeD2cXUbYUeLRKaMR0JQDuy
2tvcTQH59uWNFSMWx+rPs40CXCc69hRr/JOK/jZR5UPXNYNhvx0gDnnD3uAbDuyy
fJHUyolQ3u7+j9Cu5OBo91CPJ+h6L4bqOlNM5/QjteP64G3ltS/sJAea/FB8L4P+
3R2uKi2gAEGBr6wbSKEuclel6umESvF2+3hOd5wpo/uk1kGqbaBM3maDQVWuM9Uc
EaouY66ZqwgDXi6E0aG2OeOCWKHycyCFCeszP9mGkKHvDuFV1VVz3xF8vrUqsMFk
6dN1ihphKsSdrgkOf9Mz79EE7Y2OVeS5u3wJFaBl3hZlJsoBKnLZ0XqFCyr6wMU+
7j3dw7P8vFOR6YoX0l2aniOkIp3CVsMMMo4QiOvdZhkfn0ztYBn0PVObVLwtNCN7
Td3v0hvYHiZpPl03o9dMA7FPleF0q5W0yjx5pCq/t2lA5QUz7ouJpnP1V0TNhOIq
mwrFKapII/ljbs5LgjLOymLZhrHBjiT21lTYFF3i20mrNv54Ozh66VvqqrfeHh6N
tBCAxAsZPcgK6iZJjsCGhdcwpYVwoFS9ImOIEBhSOsKEZqkTlxXyJA+jsrJBASL0
dLwzCSKM8fM/SjhGpqMIY3G05EJXqX9FRdyJKajxEBWtFk5UsrFODY+X3X/L4xMD
OR9cUCV2yqnHhDgyixwibY2yE6MosMA/YcsH+6aaMtcDTnvVbDsf73sOskYqpDj6
Zj8U8lu49hWj68c48xGbGAdJb4ITz7/JTyjf0s8ESSv+SiqesFOqBtFr4xzysBxA
PtzpuUnNJkBGrUbS0Kqqb+VtS7gfkNp0oe9TdaqEk5OPl4dk6I1v3DiERHjM8gQn
SAF7p/7BGkSJ9FJvHf1Rfhk3z4KUYsjWljNqNrFPa74vrhPev0N197Q10mKul46B
OKxD5sDel4WMd6Hac4OF0wWm5MKMA3Pm9U/3hrf+DYY73bJsXF6SBNcj58ld8iWp
H+7SCwHK8mWNg0rlOvwlR7gA/gLEcKbsD3r/+oKZp6UHcwrVksFxjOuC5RLWJkRf
j/+w8o1/aEgMv0m/U4EEzPpO2HdjNBUzGOvxrOP53GQL0JZI7nFRFWkN2sAoayLB
TT7krLZQZyUb6be+4A/Z+aN1r/l6enjnEQo57w9niBnqQWCTaTIlScBWL8Tmq/nE
x0ijPODKo+Q8g4S2BFOBucbG+vXdAvfm0pjUF53MDt9bHnJQ2RNTDy5P3DaSA9hL
JUW0F4hif47qsyLCWe2wcQC1SDP3+5EhUIc5pCXBLlBlsSKcZU7Saq9idfk3s3Gk
AWSiEqj2JCNL1+3ATVK7v6ClKGr4oqyHQtjHXVqO6jlhFIn6y6g7TvC6rZ6dArU0
EEkJTxXpygun39hMnl0/OiXH/BK/9w3x50Ss8EkvTH/6hGUsMb3X/ebQfdCaFcME
LxzgqHZS4Gr8mvEfomuRZ8Gut/NxGqoSIRFto0knL4nrLx4DfziIA/oKjBVMT3jf
GnocfCYm6IgI8oa2fdETYH/0V9wrDd/IyOCLC7jDbz1e/Uec91Gw+ewWpDG3dLxA
voBhPC3DbGOsYJqJC27AJmqYNUPeym1CX2LImtKr4rg6WoojweikYM4+RvSY6cWn
qMfwwy9PIXyD3nl3pcOdRuyS6LkRxBMswvyqSIrnkm6kqPVgxb3KnEYaixIMww8x
QLaeteKU9AhDwzERf3wIXoYqY/4BCp3W2zNIZr5QpUzYmr5G1TBv1ck4vKed/V7q
mhmGpiO09HT2/WquItQge4Gt+u8pWovRsaWafLVN2a29kkwqj/27vbEJSA5of9TQ
VUYMsHA6V3EqeAzcSLmLOx4Zg6FE/T6d7fEUAjYxbbfJO4I3qC4MWEOUiktScn+v
E/GB1QujvoW8Bx2IWBF3BTYVzlv89U1y0KySHCb5sNirccYxcCtv7e5MvSwZ3Po1
qJufMgUCfWHybRXXNpPoOrdAUjObNdI0MV9l2v6vF+Xw1oGcg0Xuseiw82j80jNF
NglpxxWWVtRKs4ulcoLccfwpf2eJgQouvDFzABFHo9qBthGPvPaTuM2kmnjOHh4Q
yccpGhwC115KWzkCXryfB9SpJsSeEmp38X6/Ztltf+WGTOiHSG84W0/CglLqLN6S
IULvodH19iwOY5f51QJh2vlIYAN2Z8XubrXrcknfWOLP08X1+eU4yry3IBIR1Q37
fuXJkDIPkMlh1bZK2Sm0A3LFAxXPXl18Re9+rmZOpmYN3em7TY2Tzc5qxVqUEP5B
WUOlWAj2pi1deBCQFeHsPoPNqca/YHh2Htu9YAL1YLF19zvQkBEvIwvoR8cM7fmw
7iBs5ADGPF62cR0iaK7FDrAp+aZYThXyED3922FtNWHFWI526Mv1YPeibMxqSdIC
rofZpPcj8NcYNSCwc7ha3HLnqBIeK/gp5oYaGwP8Y0woxpAS7kvuX8/o5Ae1JZvk
DP7TeaMjFMzOm6AbkFt0LihyDh9ttfkKk6P4SRf5EeE/ybukbGh4M5rNX61g5lN4
ordUZ+cDoFwEesTOvP9jn1Hy4uFP3qyQuWeH2R6OgGoycc5Oak+ScKJuTslVLbIh
AgEj20lXQ0Lvu8oWTi+QeEv8z0MHlYx2fmDuA5aePj85jAAk5x3JIN/qu2stS3Su
UyC2fnJ3G3EV9LWSTe8M9D1vZ4NHtyLL+dQxml1qAwcvty54ocC07m8QN6ykiho7
eCgxg0v+y1h4iC+3zxlDc4W0pRLQWb2823uv4SaH0TqeiM8iUc4ECuNKf2RaMTch
RquwTDJaBGync0IbeE8r2rCo0C54Yj1dzKfZniEiS3xVUxOxZRMlOWP2QZnfEfpx
k+duAiqj81H3HvZa8N4UWreiRXDIAhq4JDlM1W2OOJ5w7+X4AxjZxW98a38aBVa7
arBsgdyGS5l/zHwDYCkUFcrY5gpVVh5YZRzq3e9mIrHnjkYo44MXtifXk7GDrpZ4
O1pm43ZBZoveL5CdLrQCqwPq5MzGS57AHkNuFJjQHn6/JmRp4q525sGgHrEjpWV+
kSHy3kuPvA86kUijpT1aof0DevAPqRGaqQBZE+DwSrDqIW1Dtt2Z2yXf9sKnQ3lv
GV5PZeJysH1OSUIbnwnldopxON9sf8p1pDqe+aSz+0et2CZKwPi4xwr7rm0qNPEG
UbK9xhqxdECsbvJgk3wD+Q==
//pragma protect end_data_block
//pragma protect digest_block
BlT2FS+188gA3sFfzkXsjfkxBqg=
//pragma protect end_digest_block
//pragma protect end_protected
