//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
TOb4V6+OP8WDY1kgb9Iu/mwEh3ct8MlZknQR77pgYMgR8ZT2HBDHbMB0t+Dd4Pqp
lDR8vDp2xzJP12BA2ac0OMiv9V8uNXPq88j5R/SjaJAm+BZOFGdw6YaATG0L3LWS
bPthmbLbd2nHZgXov9O9wKkBigxrJMvlPrquwCQfK62o2Vk4BZmBnnxpUN9qL6jh
YKkZXTmcGXBlgg5HaFB4YZc0YUf0Bdyul9mVynB0r4D0y+drGVrPetYu/ftx3ilx
7uugzEhIN/KH1ZdL68xSE4YkEh6oEo5GFYSfO8eYl/g3s7ybYkAHDWcS8aWC4B2p
egeiJUxnxxTgo4OpUUlxsA==
//pragma protect end_key_block
//pragma protect digest_block
FWgcg1uuwqNN0STOK3KpaRqVyQA=
//pragma protect end_digest_block
//pragma protect data_block
SPb1ebVBgv9/ZAR4WMeNe317t+y9Vo5xUSHismbz4Ek7DR1THvB9BPNHYQ0rPXlJ
ry8nngq7cJPBkmrIG3YG7t7AFKLxVGiPadx2FtgIC5upR9MJ8DnM3RMLc1qZJnw7
iaUq+mMNHgCRyfvtXJjjlrrr38l0MItm5sK6pN8vV+5B0yVie6XIerk81sB80Y1b
PrcZfxKkUyRgQx4/2ftsoTy6LScXPObZAUOsLwcbeXfE6YJc/zE7DIDuHmMhFoxT
mkNa7RbWPcno8XVtd83O1dmab9OVnmYulfZzf+uYxNTs9GyQxorPX6WY+Luy8Jrc
snjwIRAy7zfu83rbsIgotgRnNM+7trAMC0cHeDISjO/SGJaMQDzwhr9iyWIDztJ3
tmJmU//xyDSM0IBQ5vRqjIPq3f8wcltikSnd2DjtFjg9zFGau74k1N22bXCny1NC
vDM7P8iikQfuBjv1Z+NkuRSrW92OrC1XUjCrd4LfJpoJx6WZL2G6A7UujXyzEsDj
JAKCCqJ66WbqbrxDdj9SnAVZzmKiEwc3LHoj8u/GvgLW4er+K31PvVl7yDEhndxF
9wThOS6KeKOEBRYrQb7r7fAUXJmhk/mYvOcb/l1mLpW1IIIBiYDITdUSOOcMU+Jf
A8jH69Zj3duGvZoyKxXFz5CcPFyn/r1QE+NAglehGO24yOov3e+kxurWozLr0eVU
omeCQHfmLg5u0JbDghcptgMicQQ85KifFdWSX1c8MbrwG3TlTQGeJnVRHNvcFhlO
kh1Ld8EZQ25ztp22jReb7CLINum7375GMJeuatFkXWd75tPJZ+4dkD/mqQcr6ylH
0xOAEmxI0hhH6+8eemmK99HrOCwY6Nj6ia7PR+uIGMhYECeyW6HU/yNHFj537RYg
3b/ALVpU7rEtOvcFm1QVUsmS71q0V35d7e6u3vs25KkfVfr9pA1pjI5KiHrOS4iC
AjNQhZD7NcaMqgrwpzYM0jpQkN2iJasz4X1T/Vb618h831aVO64/+6YTJvP8ZCLK
9PlQQAHfh1UN6SFOw77PgJUMN53SN3bnFh08q7rxTGF8hzuLXeR3Ro8LFzwIE/sE
8D3EzIOJNVdk+PyB2EavG0yxu3GjnlHJWHUHCNWVESj13boV3FnjkI45pM1lfSio
7tu4SZFEVv8NdH/QUdxfWUafXoDAz9VUkt5Dv61qdtxB94JO9V815U6x/ZgA0fyO
tm8iTMfgp2h+fE+UjDj90my7hZUCb0VcHHVL+oxyW3a4tYuLx8Wp+Yx7epIAIwKU
HVRswE1ATZVkZf84iXG/gGKPQXTbuQHOcoYIGeUmTOQLG3R44mUEHeMy4tHBmmkJ
hrEVbhb3Af0lQTkwENZE1WDqpTqM7Cs44BayJbuKNCNt4J5FqZqr8664uhbxR2I7
aBI5l26k6INj+qRHcLILqwPxo+3gp7lr6Zq88IP10LaZw8RSLp5eX0+9Vx3x9YC2
lJTEwZaWmyE4wNQgOEr3f8khmkbO9ECXTkXoYlZBoniaD0ytZH5gPhsIUqYK+avH
mU1hhGp8btGcypNrYaola8uUdI8+15KoAhMuAtRcXnIF3E41tq2VUK0eDovjO6lY
prOwarQuMK9QPvHXkBIkIK4nKan2ybLRaXQV2CIx7DVzMvJSAI0kqkxn2FW/hn30
yJ2DckBftaXM2j+eamtTLevTunR9kyF5yNILruMUIVRNuY+/INYZ2WLSJK6s7cHS
YMZMIJWpSYtAyOhGBpfendhdrztZxk6oqwb4XHW/WVDokqRsm1ls8Lb98zgc93/b
u2wqUMWVer3rYbbET1bbJPkA1h8OVEIgAYdngmaoJviXupZO8K0iCI3K3TaXdL2U
/DXMaYeziS5t7yyR6zP3rYg2sICNsvjx60lzjAzmaSYYO07I2Ju60nu5gqoiNyhM
neVzMT6nTE4SenSSO9oXrrfwMFmZoN5rsvmYC7fZ7m28acMfDMmMd9XsuDWNNLkK
lR/q67EGN/D3aeztWKw8+UcbsWYXPZcx3JpexjyuvUcmvRTQlO6CZ7bT11/VX8jD
zyjp4SoVqSL4XZSfUcxSOrsKtYCofdfUPN3R7eET7diC7/ZfGaBGEei4cXHrfx1N
Z0GxQ98kH6vEMAuR71HTkRAHx76Nc/W2h1qw51xitsYC0Gqx/Js+BA+ua24ShoeE
XVPGbI69krEuOhzdMoR3oN1p+rw4Pky3vLM38zoAr4x8oX1Ly+vXPdwTmCYiGcng
XzV+a5ALg8VUoIx8BnZ4Ue4ogKZMIEqRAMmgm1wrgLNnzEHHQczhwZFUaCwvKrJE
yoiZORVot3SlNrfMra2umkNctYKg+eAo21TMQ45cW3k9lhicKRU5RH5mGBObhqMr
eoABWAPT61xPCFuUFMgxEA4xjNKNxc2xF2tiext/Nx9qW89/lqZOIzhtAy7Hv522
YF1eNuRJFpqGpgvrs9myKB+4YiTNxS59EWqyQ2d66LwaNj2TEzsKQHL6XYcOqUGA
0oOmTOnQEQnq+GiZPO3s2EVGmOFWts44NMcKLK4xnVlwXRBfHDSHdUFoja+6ziXo
gVo/tiD8/A1I9M+PdQmu6Z2z7bu7G+hYH75M7dSwJ0a/Xb6RLe0CO1wjEOsOYULd
8b0AIkgG7IY14S8vqrXsHBqfV1yX192O0R44QJKN2nq5tmeS140a721KQHkl59MS
mUKvAX23bVuF1iGhUJ7AIX1reRZlzRG0CtW61tj0sE705W1Q50UzTZg6557r8U7C
N4Ve9qoVLE5x47J5lXlmH5/IfZJ4R2nKS3ddr0WY8pS9GUhgVphoIjfjqWrUNxSZ
kBBA/wYXg3xE+fhXwCg0Q+8+ZH2bIgGGCS5bO/VT1ap5wHgfk17EYyA8qHMns3+j
JJ0hUdL6Bw3nmoS2FP+FjMqT/O1snk7verwamM1GhSQFCCeK6lj1JYbeuPhwRzL2
c79T77NG0vuEPrUShl7cqduyUjfWjOoAZiu2XWtB3IktmuKmu7lf9b+txejhIbCZ
FEdQzPty+jptoO12jy7WJjIutb+4f5gS/m3o9tK26Z2gndO7DDHdlsNDAlxgkc8+
JWISx/JHelFcKa2a4vt/nat3vTgdiZQJnDjhxe6PK7Zi8bA8VYbzj8sAo1EH4pUo
MRDNeU5CuxXVA8wrTN/chv3KLDiQiAiKmwssprBTc8fJHhLP3Ux8KgztapbOFfn7
t9+4Kt1r/j8yaeVbtb1i4sQcRqQx8R5pJ9gvdpdUPo+2bxwybw7gcxQEp6Uu/NFf
wlkK9nfH+Ze3lSLSZXDTM9X45cVyzMLgOyOaPMHq6j7CxC3/NqpicGLCnW/UpWA6
q7KZ7/WsJORlkiSrz7Ujxx5HV5OTq139rG2PRVfQ6+Tj9uJfI20W41JQAECvaIVy
XmN4tYMIhAZnrgTkKjI+7HM1f3gxC0LLGi+CWwXb6VR176L3aMEFszI8I1Z/WKHE
DidCJ0qTdtLZXmQdEyQFvAaBRvf9p6+WZhFkvuWSClBa/ubmQaUChZg88Ruc2FoQ
V9r6jdIdfBvEAAqWZraeh/X2HSoqBrQrmpXxAVw6lTyw+qMlT9isFDfi46Y0irHL
+zYPfBtOpmM+QhT8rIWCpB2csjkDuqxKU+Zs6ey++QIepSpXdDCavZULjuzXUQr3
DRHSc93ypd4q8uxn6XMMNrYblyMUKajn4eU+T14hz0W+rcF3LKiwYUzsTM5f2fY3
WyVRd5MTD8RheUKq4luKKDIubtfIP1fTwk26AFz7/unpBUEJ2GJzRnssjFPtEqxP
aU2NGDE3bRKQQGR1cIfJ0+Xl8+bFENTXbH2Mp9ZiXmCFGjzCFd4ChaWBm/94alGX
Wavlq9grLTjVpNGh5pjBfl9p6fG2wp81HeAsqlKMBuGvue6NvJLmy4vBHNkNTkEV
KdfrNwQM6lfWZLw1XWluhXvdPFSlUhmEsbTVeM7zIFDuV3snqZEdgA7salfp1/JW
JHsbvjc+ntoeYj0A5dvPeyDusiiJd43TuLr7kGpo2A6uI5ORRqV2CcL/Nt+lKNPr
vLkuTbU6H9EKD2VhzjLDXc2gazbsZpJA072a7ms7Z6neiIIsPrZpxK3KGOlwAe84
YpeIvkxd4cSK/w6OCwU37UVqxWb4cTDbBmng/j8KdPFwIegsnme08Z0tkhEnsfhW
I+VdL3YsDYujKheCQQX4Fg0LJVKY4HwJJu4DdorbtrzBJ8xVL0ZoYBiIa3uEn+5/
U20LDj8WB7gJDmxXHKqEfZ4fkpMhU3s2xLbkaKAleiUxmfDs1zMTWuRZjzeljuVt
TM6gP/Znk0+FWRSNO1wjFPrOnJjmsbTt7oPNlKZejjk45sosAfdUPmnJd2i6SLcJ
UMgIYP6KePHLSOJ30tqxdfBO5gISEgLpUQj21i4NiAir5nRaVG+yG7ke6ExePlEk
S8caiUbBrf6NYWmTn2fQuOS4R8PgW4zk+DDAotApa1lU4clce1UfyrEUBCFYKis8
YILjDB/OrVzeZiuaTiuJeRyL722MPlsoAckXAR9J/R6oK7/E5Wk83S2M1f9Xnlyg
CXscCV5D9LxyfFzxUk7y31e2XWcwB4qOQNQEpqPCcfjkIGNblpQOLSE3fFDJ3cyV
jppjs/jVNs4vdcAr8qNyJoQfeYbPh2uaegFpciuRqH2RN5RDY6DXfeaVzwjg3RNH
dgzPbwXos/4qzyK5yM9gZ+0Rcr6qdPKOkNSpPUvlAhNswwaE7nF+4wAoVOWQ3f+h
UFOaKCsoESI/W832lTuH5faLyngBI10YlYmJ4wSPApCh7HOZBn4K1PFC82RZKM/X
gdJ4we/kKefsVFyFgWV+F+H2T6InbNCwMzSbck7pvlQ4ormpRw3+rl2A6br6jHhe
dPejxcmbAxuU/8ZrZfOn6fWtRXBOxO4eKNAZt5+k4rrvRACc/CeRlLy1DwqoqrQ/
LvwfT5bqp6RvYi7H9GivKM2W1Lr/FBn4vcKxYD5dH/ZrWxViXR8e5IIz1HMelLZR
cMpNM1FwzAK/ekZKjpkffySSvcCHY00kmjD1D5lFSJ6pmi7NNKKJoTcmNlN0AqgU
iou/pksMXWlz22lW9RxZTs2PYs19N93xUjcohLco8hp4H+VJRUwMfLPpCDTM9UOZ
YVpruUTgt7tHJQYeTAtujD3lqAafus3N79N+c0dAp5DMED6sPzHnEB5olRMgvljr
Sc1XnQb8m5ko94WzW5Dizk5ueya+1St9VgSUQ3u/S4GbMyexKNHVQfAFjkJfgOue
kY757TICA2BBgVKZnqpdwSv+rSjizbzztWdKM0///cYQr3GbZUThy6WB2x8hQj0k
ACZEk1atXQAu4FYfVPypRHsb9T0kbir5kjmnLbf0v1Rpfx4GpUSVo5IQBaCMtRQs
BWMeDr94ShxP8UQ1jULVycgf6MQBac19/gPvTeKZIkiSBrQoP+BAky+QyHdjDMeX
lPftA9KtxeoQkm7PcxG9h+hO+X9rTRFPU1SOwDbXJho/9vWdVpdQKytlxgdpVWv8
LrDvvDk1Z4UHhBevfCSIFtKoBcs4gSkx3/D97hCJxw3VNOJPwDeryRsJIOu97QAo
NqC9Lk1+JE1Vu3rH3OS1AkrJjOm5WOzkqW38ErsUnDEMmv3uhAA77flxF+MFw1Sd
zb8+lRHprVrFlWoT0Rz+WOs9obbXsOuCYTdRdgjtFcurk6cxx/GjparXGXNch604
9/o/9RsYTG6Vqk2QGLs3O8tWAuwPZf5ZbkGtWwo9FTlKk1DohOo5sjO9KsjShV9K
tWvCyAfZWt/xvst/EJxU00faZekVBTlsVMMyxBKPRVkA4XpK7NWMcYI9WMZiKnUQ
M0dkkiQKwhxxJeymCyfN/zjPeW2jMJhvp/0ECiALALTeEPLDLG4eRexTAz4SmjI/
SU7GgOkmlhbuEWaNl3/DL7yceVYjmJ0s7wRSFG1ZKr/Puoh93SZgNpRCGUaOtdLI
yme176qHwhWlLmuVFOkfksBYsjZtBQdeXaXvXhQNZqe5IwN9CU7/hb9x51QohPKM
iK036D4Ic/AhqBJH0vV+fXjAySVVFk2SkooaM+kAqy0rDR5crLl+Xmuv59Uuv4PF
ent5/gkWi2sajmUXZNZla09VwO+lZni51gyPalhfpzyd3J2vf3aEFRCOleTKv3cH
36KP2z67uI1UyvhQUn0RNqwnu76l9y2pMCb2KR96Mm8O+l1W+c6aK1wjJxlrW0jT
PdeI/h9LxSdXKu3bm9fzEFGSsGU4x7wG88PV3mbT07+wF+7SWZSaNwpmnUD7f89U
DXHwVXI1zLk9MhstqOGN+yYAQKmDqiUpSEEjW4w0Nceezd96O9hLYobFEn7vqFQi
ChsSpz9YFwDj7ilDqBr5CT7qENoyv8MAPCseIlXskNM85EIu/76w5pQbvkD6foRK
ZILFzjRVs3qZpcvyd9lk60WEntJJWNrFuy8gVef3hztcf5KBPzHNJ0+BY97yYHne
N0ECUqjRSQUHAMnxrf9v68e2oBmmfEHa+n7wfozsn49pP5WK3AfvFeOjv4j0913Q
UuBhOUor/jeSwUHMRbMfWGoYN0vsZHCVuoSTbdXRbTRMXrAk+DslOU8QmOBFTpMD
xyq8bGuTLaUYaZcs6Y0eg88Ig+zMLU3z/11xEp9ZCyGZzkNv/qFF9Vu5WJLD+t5r
wIAi2QiJ0WrnTRrfzTYlKztGh5+ohdhKfJDc8d2h3RaJiNSX7zK38glcAGQe5CdA
9SjjYJX8znUbrs8NBHNHxESmUinSX2lFpkwr4ECd+mQJE9XVakNs2FuTcy3p5B99
911dxClb5rnXix0MRDuaPYd057F7+PmWP+9ENaV90iLYGTGfTxMJFP4glyPpmwON
I1+3drmgSC/7W774zsl+kagaGZ0SKkxuSogNiCM0IkVna3uRo85KaYv/0+tFvOEv
+p5C79yW1kLC7tnU3us8bcyTrto6gpm/QauhJpY+3+d3OPvEMmzXe/TW0LWuNjbD
eUUbU3I8SsHSWxlYkrdwwZIN9e9HCbSUJr8R25I861iSxj9whFC1cZ+iVDOztxh6
yxvsFTfR09TeAnWVW1Gqd42oF8YtvCHMRbOMcDHLdDxml8Q732H7WAQnqVG/Hf70
YXkMGorMgv295clnaNHYg8zqobnGgjNrpn2X9q8S+k/2dIPdRetNRqBgl4mwcqAa
dFBRs647tkxLIugUHEQT6ANKQpLe5xpYqZmtiVxy1YXqW40oTzkXLKn4sNUubEfm
DomTCm7/5jgqVdqk4Uo1Fe2lHdpYro9sXWHiCaEsJKukIlBn4zjib7FNz1wyB5Sl
jRnfqJq3AUpkDrMWqw3SAaxrHaMNcGHi8X7WHXlvGD29GjMPdf/7H3glVTujv5F7
g9HhX38wuvdlqGPOWBnjYNmykyY5P2DBjObvo9C0Gi5KhgZU08O9QoGk+L23BAjl
DFx1OrmvN2SL56Dc4xDn7naHvf1YoENQ85j7dThLUGAV511YS3pHaxmRCqGwmmIu
T9xSKcNUM6ktldG+BV5YZyJhl1T2Lv3VVAt2G9FzVH0nQZU5Z7Dx5zqyrGp/75kQ
xSrknwvWnx09pfPf2YsTrGP+ChJZKWuNRytnUhvWiJeF6gnALp9RXBDyMER3nf8l
6cIkhCXrOQEPWpBcm+f6WCJlZ8940iyAClytFqKH3UR9vYSdjWiJNT9Dwi31s7eq
hRl1zzUw/r4SL1P0IdSG9PcMxFVGEQ8u5R8xJw1YWWQWbzm/8XrS/N4vPUEhkK7b
XFEpFaCUb4bqoZbwlyxwTXYA59yv8cek9pVoB0Y2WfiOT9+u6auFZLif/siP8x1v
L3MSJdPqClL3jBoZwCtZL2dNqTTXi1iVxysdbA2TwkXcyFUp6DIe3Rm/X5rt/Dmg
1EgOOWEN1ls9Qk5sBvIwqMD07agnsNu6+Xk35Qr4TqBBtKnAMJAzdLlREaWZhUyt
wOsY2mQaPEUzA/7D/alEit1k+c0fTNzFSH8U+UGWFjx/kWFpQ1O6GUUgjv5AIfx9
wgc6yPyrBR0fXqpspit8mIgoAJRfJMSTjhy7Jk947JZQrv5pJHry/JhkuD892t3i
UcIIIBEjpRVvBGFDfFaMXU81EDUpMsv9vzqwKd/E8GHd8gfm9eyb/yIw2ALw8l+A
qXpd1//znkz6PuXf/MAwlbdm+EITXMgKdFHx8ymf9ZEeRSipFRfcRIuJGX6WhY5C
NauV1QGhK0TXY7PS1lsMk5A7n1mw5HF8ZZlYXnD8CQ2W7PxBntPD/V3JFmWJ5opq
DrlEsz8kDymHjLBdpH5e8djgpL2ckVtmOfaDcAVnMn7mpOT94HirPFjRqyyQtoTB
EUBP7Dw8nw46J0S68ptB1/KTwSKt5hC+wkmJCSMWKEvivudhGcX/ND5iUX48R8Sa
zd2X8AeSwkdQe2QoRE4WE1gFcRsLohMlwtRrf0ZOrWPD/hjn7c1pSKN3ntGAIOV3
tut8q1sWcXlAkz9OcUW1CBx9ZrsNwkhQcHWhL5nCQws5OmkIPmYf5S8LiUKiF85H
xB57amX6z2O9Uv1iNwaadazNn+URmP89Xcg0IqqPRY7iT/28pJRJNkAcbAJuUtUA
9iBZ1mBrevyeQQOneCIEe1nXzIf/gX3Vx3ryJ6P1M1/mX/Xu1fBK7AyK3dyy7RO2
ApXH6Vfr//lKOJZnBEqJo+UHyKcExTtFgXIgPGGYenD//iR8cUzvzG/Mw5Y4+u8O
kZ3MaDY8fZISjGFBUmjVezjULEWg0QdKrbGD3+djHK2rjCJ3EhmiTncDtlELQZGt
t4oWTwdHgsEhY6rU1liHVYk9lAJrE2wmVHGZVPAi6Vd9w4tc/ggjTZgNbhUowrb/
FyuxmZjdSQLcuoL4L9Lwwa0RzDdM6ubtWkkyvfPBPUVVOfHW+Ef3kv6XXTfTt0ht
vwnZBa0I3qN7kzXXhJAD9nMBXtRtEFhThR9P4Pg0LBBo/w8IzpKvffwBKO2XI4oB
43+rgdOreEJ2nBzvDHKRPKexVf7uL4Brzk01LOclE16GWWm2fELedCNtLnHRNGeW
jsx9l4N2D0DPzt34vVollmb0fmJ2zllK4d8/YyBayDUhGDS9TEuGUOR2OsBdCFWY
pnLUz7R+NZ8qZ4ct3DgosPLoGP+rKfwXdVy9Irs2tm0WO28v5/7UJbGOts/uHcsE
QUUojxghUdJwfpTqSv3jb2lPD7GJdb2tyU5Pt6ZAavyqwJvVy0EUoAYgn2r6WD0O
pSDe4VxiDfuO6lByBa9q3PWOVuSszvnkZvo/hK+eghK675RmlOGzVLXH2+UCfirH
/ynix7M1hTwlkfki/+i+0TAAqw90b5J5CfBDhahhmKlgddpaQyIA0ecCXJSXaCUV
wtqFxUY7E85ZLvsPRNzv1Pi5RXsU+IV2G3kUE4WXBL/RxSQdv4WQO8rovtlTVmgP
a5UOkUylUgWbSsqkCf8BYGWqhdFNzuKdGHtqVqiQW5UJvHNLU/birQdJ7CAOOgb2
vYervjNOFgIo+wEG+skIOqLoUVij3PVBslcsATq2+7x5cXtNSgkvfK/+L0Xto05v
c+OAFDdb70A4bKE3jFwUQ2ANe3sMEFQ5LrtCAcKYfkzfGvKpGuB2TYTOI/c/0Sxm
q1R/st742t8UDvwVghejh07hn0MXEitrOYjCyLQizrP+3a3YMBlvDLdLNhzLchh2
QV7UhlZZNVEGK6RfyB0NLy2SylfkuXzdrE/AMDg0SiMB775KJ2fvnRuN134MIjuq
e4IB/0oMSCYPA8JMhRqXe26mEGjZa9FtWRZz1xUzFgzS/WEKzn5YgHbDkhEg1smY
779tJKA2ogHIHj5v6YDG6bjnMvxj6V1EV6gwpgfSIED8J5/eVNkxEhkh2LKFmtLf
+pAKAqkzPFa7CVJVmDmCHlRqHQdtNw5jWG3UjM245qslSe8P+oLjmep1gvaKz0f8
iaQ1wBs24ULHEvNTo/RaglNaMfVnAsIVXxvEzBgtuU7kD7YL0FoOVLG7u8MHk9WD
t8kwy5fhHXecaMiDIVzPJVitG8/k7qY4HAKXyC81y6O4+sMhuULEHUeDoHp2n53N
z8uRcwxgoDIFtGL7dNf8LdusK+f8ky2VWOzvO/K1uNBEg1lKSwXlQftcpuiMNoMn
3ywgf5TCR4+yWrfzLYm1Dumhpz81L9jNM+x3HemJVaNWBm1QVCcOc1AtIPSgW9V9
kS6jJb+k2Py84BQ2z92mckla4Z4AEBhARMEWEthgMn+5hv++AsNRsx4D1Nhj68hj
OGTq2C93QJ6OVvGVUisMyxDpvqu8pYZaw0E6fZP2cy7XuTUW7Q5GVA3ok64tH/5o
6Tm0gMS81p3ZK6aqGytyl/G/0lRkibt8m4Cs5XRZeCxBFAELLAE3bsMku38HNUcT
mykEIgZFWiCRxOS0qorTA7tRtIvYY9ikXcTYnPpj6A1dGB7CzkFYIduXhvtD08nY
rG/E52G2XPKrq4XSibtjsxy6Z37plZvktZhOhirGJAHvVCmSpb1xLuD+j9Y4XY79
3RICRNWMoo4M5DvZCxE2bmNKGq5rdUMlQnToiZpm9qevh/KqGuV9CrrZQINBvLKH
xhfuppaPupQQh37PbeqgBnzv4FGIZt+yH9aYSFP3hfbbsatbE8ggf6JOmZlX88cO
V22lIiMCjyWcuciMRnHsZro7RT6atruccFXWM+PWlxHdc0Qb1y2Kjfx6K3dBbJpE
pqUO31d0ARxoSfsnmIAou8HostnSnIH8JIyd1cQX0rV1j8VTwZ/orIv81+GoL5Dv
8SHtu9pZ2yUVqjrMDJonEGOGYrNXXMDOnibXgtUY69Sk+qWtwkWX2fjEKgnKWGH1
KW64qoTMOPhPBanKEhikWnCYk3DezP4gkgdUG2oN5TL6fKbStbTVBSEnMOMcs0Hh
GfWfEV3yKSqdOFIxlce837MR+4STPLzKrHIStmYBU7DI7JsPMQv1ETqv2I0kqOLj
vkT7v+cCGmva4DyQNx02yLWmAKGVjLSLTno39qnbvpPI1VzYHC2XPRG7Uwd4U8g9
mgri30pgZJ15fpSB7uamlWRHjTlTWE6udz5llKKIq3AXKrxxUtXuqQrdEnPRyS4N
HbOIOiJ1eRzSK8FZOgZz5u3l6OBFWwh9cMGss0307vcWPyoA5zIaX/bHSHRsqiiy
l1El7W42vRAOWKUsc7YrrHaNorRH5JA8Wb4wLCFa1HzZ7FJNv5hbajbOBs1OLpWP
turQFizr8hGDJ1JPNBRIx3zGmaMzBPZHupcW1DOU5vNDQD414KXr6Ge+XseQdBJN
K0W3MitCjaokLv2zWDfvRLO+Dn1Cyh3ijIDYRCIl45orVTq56ey3F4nQMhNX/9rf
jxwx9+Bj8dqjR43StWjygTqifXbYu45cUY+NY3OQfbOLwh0zeMpIZO2pbmwlUZkc
VlNxs6kJAZXS7wXD8ta7oQCPu0JpHqV4MiG4WA2pHsCSAjawYjJWB134Pqu46fiQ
3pbzAOFgy80gyx+fX8PbCr0s7Axf60tg0QiJUWTtkCP+vdGXDcN287TbmxKpKigh
2tIcZ7a7rQau1+uQJ0+GrR67xrCD7W5OAMLfLXttbRklvrGujXxmDW+s/oLYwrP7
EHG50rox3ttoLvUCUGQVVIG+GVto/WsS9cHnaHxTS7Bz7APBOtPWZMM2Okv4Ly83
3mxDkxJvUi+kxitof3LR5daan3u5EQJg/s3xmHBoAgT8zEBX0xJDX4Dc2AKeGC5P
rcGELaNZHixnP8yS1cM3u1SeOgWT4vK3p8ZCO0UapI1pwiY/SxeswumbfvaOjsJ2
878zBSVHm93CagSbpOoZBnVJM5AvYFpaLIAeaJ4GAn6MBKMrYsimRrA2HHyPmdUB
nmorn0AvMO7A94JSZGiJLZ3M/gCFhhEeWXL/HjgbyAtJVFabSZiuVxZzMc/NwEzh
RrWQ/CtEtBlKIIBxniw5hkXmj2m6VrBqcW9mT/u77Nnapew4hQ5rxLtcSDMMRw93
oiqDoWCsXutWOknKIa8xxcEs5CG+sz3Fx15tqxCN6Hrwl7DwUx7Rw1Sd/l903ung
w6AhDCVjbqcCDS5+RVaWBzjS2CczAFp1pcWDcTw0sYL281vE+L1+Q4J6FyZ9NMuZ
cBKHhp6gy5uhhSpKMCOJblx/PrBfkXeHkW0IU9b0JODbFWYt7iconRJxfT/NHZo4
Vm9JbKyrRpgOQNzHTS+WVvAy+EgIY67nLo4M5hEDZPRvpdZxqK6M3PwOtYLC5bXj
EQ6PjaIKhngl9a6BpVabEkGgBKq2ghz75OGJG4WEtnpwGNltk5bmTLy2eJ64rSKE
XJzX3UhKV9zT4bTqkZQ12NdeYG56kDY0h98hKDRqtruhnOsTnmVj4Y2+Ha31ezQi
KPuibYrB6oH9W8PvcgPzaisc4LtlHtnKu3xvQ0AayJ9xG0EwW0gScM5i8gH0jKkX
AyRh5mDit2nnpAcIJ8hvh0a+AvYs1ilUVaYxYcWN6MB+AD8cnEhWXI84UebEjkZY
+qphEFV9Fsc+iuVNu9bzKNTltmPupvkiamJNdxofYZg1pGM+Fhk+finT3gVGXfWA
din7EGcxIQNL2qfoyuMIthhp8QgrVAjWQwA6hgjkR22O7dZD0Dzw1njO9Sy+2+f9
cvtfbw1g1H2dosiNa8w3f4gLnBMurlQRMS1fvvCGzhnYfZfo7HCG8vPO6Vu8IVuG
PwVeKVyms5StAMacDghHz7LsOKT/23iLvCfdsn5eKgcGC2LlYhQsq1wKuquVai9B
bmeczVrL8FO/VTBlupTXBJgS7XYxzM1LciGFKDLh5watd6iLg/C7vbmvl6KZOS1j
DiqOpbQeIc+K6X9RWsFrtofs1NnufblCUILle7rpD5R/DsuX6CW/n4MlcKmYGSJo
ben4yGv6icZh+qd0eg0+JVCRvVvYsGIMfa7GLWPdCgHfsSx7a8DjoTwJzObYQX86
hKQsKSYRiL4wXueoRAHbVk1rVKg587SpqxuMViwUMKVSEXUNXF837scWQmorvgFu
k0uik0obKVaXAYu/lwYuq8SkYtQUr2ZvLYIyKglSvIFRiVLV0QVu20RvTN79q20g
u4Qaed15AOQxx/3eQLea1w1JtdEE33HzrwxYfN56Oe8aRBg+pESw2lz58jkqvjVP
mkyBNqUnXV0/OES3ZL13ptTP7ivR79S+6AQU9hnt+jSX/dvHtLRSCzyVHCFu8/rP
9xlGlO6y+MIdaP0HTxijppD90GpVHxGBNd7OlXXRTzp2kQSpdUV2cgTko8Y3gsZm
RG5gp3LIGTdcPICr17dwxJWq/oGBI7xo1cTp1lLxcZYZAnRFD7HO9N1cFfE7Gm+f
br2p5pUjtIYUmGVH4xXAoC21j3itLExTkU5itrkTg5x7HWQR6pvJAfzE9o3W8dEh
LefYMZD+ySmnaBzxqAzrkK3TdDruifKUtB6Fvd3V2vbZ2ASWXB9wnXZEj5sycyxz
icRsWiqpLLvIftiCxrSncY9Usmu/cyWw7lWKiKtdAOEHJPooFEjHwm4wzeQjxiwj
2x8gAV5tlAOUTrTRoyvk3o1JQ2FN2bHAciwpC3mMV8mnyocBY9rLypInvig7CVtv
jLRLIO8vDXvGlGUDuARER0W952A1seFbThtBBvpnxp4Gw3p2h/eJuaGdGZKSDGZB
NsOODAwl+XVkl4pDnJ/bfHBVu/UYlY2LYZPCVyflcT5j7Bbdnt3YIPvD1OYFH+Wn
lThr69Zfmdzjgnij10QzB9an869vmvut+uyzA4vOpPplkgU3sjutZncZGcv8Mo/r
9sQW4jYKFDR7JT4SsQC48RGY2Y865BDGMcEDNGvaEIEDNTM69FPGZU9x7IbBuw6s
VSqF4NdQvrT5on75uOQpb1krOTpMM893HeilAngQysKageJvqKOHoty3P8TZgyn+
GzDREz/j8WbbTpQALeeSPmbHPtXYXohtf3h4o/yUltrC21RqaM9BhQmKroX8CFBS
VuLUSwuoreUVWX6z6OhYWFV5p6Tq5GPsnczrxs+8fW4JkRJtpH5cfE/nt8sRzSaj
tBpVy5wKM+eendDRRVToUjmcotguYSKkXcj9XklBXcnqcn4q5VUM+3NEZQP/AShN
QRKVTX0yTjQWbaFVwkXKSoY6BY3+m9hpFGvSSlYRerWTSxGcRmFhlTIikx2S+8YL
zlYROATPMvI5/Kbv8Xhr4XmfAI3BbMib6hOgnkwoo+jU8otUocvux6skzhwN6OCi
lsaXjtX2w2m8TNYI/ZDjHldNuiXPCStGu6SznVDf0HGpnZ8nap5SIaPf4rA9dEmm
re4krSibdD9oDCLo1azla5QRh5efhCKFRuChinIMBuG8yQDF1Q9DNvMh6bMw4yAD
1lzMYQg5w2JgkJD7X5rXnhZVa6KDS7w0w+bmKnMEoAtVP/cU8e71AU7lIP/XCHUC
D191xNi+ly4xjGtSQpfQRi223aTlx7WxewzMMgoDo4m1T/NwxzISYfpM6SyrJPr2
yFWA2P3oCl0FsW+N4V7KTB9Fr+zeMnK7t6mG02mfMTICMiRPUyDeg8hPCPsDYqBY
UDCPDvouublELAVhiqSXCUnY5SJMJJaEI3eCxjTgPQsZGtRbN0Xq2/nlCeJh4/xF
QryxP3kdKihQtV7GekrxnIYMcvcjguR3ZjoX8/GOvwE3l/eqUyDku9rkxbAnoEIC
usbfZPcj4CcnHtyTdYEpJLXTSB4yGCuw/P8a5FJD0EIXHr1uF0QT9IloJq3Z2D8U
tUys+TC8someIsxepi9ZMqUSYvDn5gAgN1os9IjghBUCR9ufFT3m1WAZ9nxbz05l
csS2vfa1nXZq0oDDmzvRABOcmCOXFgW5aZZxL/oTHriqP3kt4woU1hXNA21WeRFf
yjpBXP0IPzEDWpgczkzN6wsP9hFxoN1V6yuXj4sRe8E5e6l+kU4eFrdhgyRYXyHL
BqLRO9dddjchpzABEvBLWLahB9d8J30lZGIfk2WTyYHmrLpe7Ob7QmwLojtHSLZP
DxUcnEjb9eCAdaQZEV3iHcttGmheoZWFM2H3g3QKidvkAT/CSkJxUTsJjfN90Peb
0leE1F+Ge16Op4x8vbWpVOfxlB/Yy9NA5ywoXnUOYPJFzAXR1CAndtWZgSL/Hd84
OXaK+vZIRZKVc4bTPn2jJHERmcvUTuYJFoCLtVdi3MXCp57GdkZmOwZya2j8K0Pv
H87lCfpzXocS0qPoYe9zHxYE6TLgmL3rLTKlOjmqitm2oNngHFDiKOYn61kXeQz+
AXSBdy8vov3y9Eqkwg5pegSIOpZ24Vyq1G8ugkZC0CXbBALPfnVyRMrQ7NiWQ7ti
3fvVYZjP6KGHio74bL2VbdQoBw7lQQb2RpP36ZNf72QKSmS0aLx2J3S0PK/JSJhi
SrV94uUAHgVUh05r+V22qf+9ZZXmXIVwrlv3JtYQFZnqgfCYvqsUm983kw6YHZ+K
gIqV+9xLsIP0Nx6O9T7p4nPEqn2kz9m7vaDDZvh1Z2liKaLJcpQ+o+qV/h+rJO3B
3TXr/yOP/N7WHkVbZjR70cUsu6nxZf/9qMCmQxpy3yN2pOsuum90RMn2tGR3d8dD
srLAUxd/SH6R/okKIBYHCR4OYE9VTbCcsTxvzSw+Ao1OohUdlXI7vtTUuHw/Riy2
JugBpC3MZ5cGkJaD0Ys9JhxcjymZjhqW7c76qy/DY0Ty+9pBuDBstai0owqaFJ4T
OI2jAEiwC21BRBQIMJc1ujDB6sLd0QGIXC6YbIFc+00ppeHecTQFuHfZnqSs/m6T
c+rQkFJToKl3vCWQWtSdvfglpDmJjwX7rSKTq7RgNQuU2f2un9d1x4gKfbpYTQYf
2ahH68NZUQtWl+dTE/T5RBXr1iQxbeAr09NYQkEFU0eQWA1D5Rasy7JB+Jj76qtN
4oIo76r1nXUj/JyVa21atbXF5I1YR/K/ANqo7HIkadx0ev0eopKa9HhM5uQmsqE8
CrvEXDQiCzK72hTWGYTPyNqHY0OH3jkdwE3ucoVem/u7ZUxDEYmqYEFb5kzRtXKq
RPcAVS3PDj6WTgjNsQcj9w2YVXTQDzUUEGg3eLuYwwrAerV9V3VTtF0H8ifOpQnL
oARuybLjVI1wxHgzWEmHRAm7Sozsjz9v4T31dRBCD/bK9kjki6ViBIUvFeAnsq3z
yY2CauvUtPJ3Yc2Gah9TnT6q1es9f0iweUdgC8bObYmuYA8F6zIvAcal6LMMF6vu
zFZOAQzBRH/6FfvQ9jayHrGaLN6m0Pe7Pw2/s5ex77Q7rD3EP2JBUjiWvrKDEzI0
FW4H6qxUVaO/llahP5220lQeAYFw0k8V5Ln8wWTH9G67ROUPXVvN4HhCTu46POJG
L7ODQstBHdi/vVlnBSV4aASLSm1ftZi2P6BaqP4JrBbaqy4UfrYxdNGCtzRejDWK
UQKoqE3rhq3x1dhb4JWvID/y74EJQwud9azO/OBvfEEp3poEEbfiKPOVdbmmrZz0
FfCRCYPeGPDms24+bQRfyx3fj8DfDTnKb80CYoJlgPiieX1/z9tEzxQZV1XihEYC
S+EKvmaYEyBgv8hD6ELFIr9XWT2j7QT7uTyhFqr9RnxtoUhna/GMGV4kalq6gD1K
2YwWYndEV4DvjTBm6KMBzW5cqRkUW8znfNBKqy6UssZvX+MzI74eU2tHvuzZqUbM
t+fH24HjCFaXsfOxDL1A9GbumYZ7wKdYwh8FMJbaA9SOZF3HPE8OQl0qpgVOUAbm
xrR5vlEDNHW+PgZpBbOchU9Gyf09gGRVB3HSaPSmxacIfWwuJC/4LHlfYrE221UA
8ANA0a8CL0aY53G9lxWDk/rCnxztG+m/olV7kPsH58MZs/wfpAltwCcoU5Zk3TXA
QL3QhSJ4UooCjnKM/JLICQIw0GjI1H6u2uZjc/wMmu9ip37Mrj8Do2HtRA2RkNQ1
gjuZedfqbxW5M+Y9OCnfvxbBbi/8z2QRuuLLrFJbUMFlPuGy6N5ClfY67Kk5eTGm
LNi5Gfm3nO1HLAnZUE7VlJdT14D4+qJD+Rbq6jsRQV85hFCRMdXfRxB5a6oakgD+
8MfibHA4YeH3dQkwAlqwCTCEQWV/9glRyTdHkxpkfW2JbmPadkUO+xjI5joDlXG5
vZbecT6clSluu7hjk4kTLcZqkUCfR7kMDTd8r9e3lWg3fSqPuRa2PfeNg3CvUOk4
pF6bkJc8hpRcmvdW1MLZKOVN6Plcy5E0e0BDWWx6M4pgkUTFJV/GCm7M753xmhwA
BqPfrVwxm6EL4n/F/Gf8rZpkCschGSI6xoNg8oKNQ1xiDW8FZEW+lHC0KV3tRRsk
//D0IXXnsZ7m16bmEQSvRpfGmls+jt3lFDTJjGa/FGWAd5Qer+gnGMUfXVfXWioR
UTcy5QiBV4ts69aKg0Z59S9d9caLJ/7J5UxAfWE5XZqEykcguznExy1kd5whJe1/
IigIZR/1kQEWKgRBjc/PDrrM8c/qd4BRtPEOEIC1GWcsM1SxnhTPYYvLDh9Om9QI
wiAUqB02dQ0h8Aejg2lLe/XzRR08dinm+r7jCmY354wsO0/8cE2Qj5cD8mTEslkj
ASw2ZYk8ymlXd9oCRpEB9K17CPXslAk8jqZB/wNeueALijwa/u3ZRBmbr4vzOoVO
xtAWu123TIbAMOudIEOg7NSq9r0gt2JiE6AV7OASaXIVxxE6cQzrSW2wBkSlK3va
1wEgWo3SHfdgsBgWxRBw/YKIs1+UBWa0DStP9QlL8qTC4+AcoqBI5aJBUxx0QD7b
/d3fah6RbuB5vJqFxk8cPaOT1iIMgeu9TQPnyO0X5XFJWm9uQlbHU1XcM5QyXBHZ
dVe7XE4bUZecSnwdpNpmNZi6oJg09J/VFoCO9hLy9l0NSYaw7EfQ2fthnsA2ytPe
SpvYdFEbuIaz95oMR3prAcAQXdXLu63/Voz+qZtIWwDbKekQtDeqfSb5iapqtw/M
jbhRzF8VaVQkDojjexjfwTnWUb8ybeb8HsRCVy2fAQpl8RFtlAth9GY5mIV2FdxU
qJVgE+Q8zJsdzcQyW8coiEb08i+1uqgecmRIdw0TzI9I9nRdBQjW/YanIAV23k5y
QR/dJcJq6hADncPur+X+6MOMdBMp865/ktHo5sD79n63+r3ay6tOiCo5/ADaE8Yj
uQdvoXt+DtvqnzLqaNbnqv+C6k3V7UyRS8hmKCujeL++TE9GEt2uPvPWdmLwkRsP
vHhHiMHEGRfcqRkk0j0WAEoZ7mkCFrSM7DptxwcX0jn0WttZkyxbgUGvuWnpakO8
HZHJ1FIaX7ILxCqpMH0yEumVXnj89oyifD/StFIhI5n7ZlLWgitLtyS28tqUt6+Y
FGpGoE76xzcJ1FmuVuEmDjIONCcFjr3QkoewvkSNvmXKFWTPSJpeN4J7jWGw8Z3N
5WqCzrWAjUtVMLznzLHdhYJ1T05bS/rdb7l9cW4x8zGRKhwGH9ZlU/9JQUJdU1rY
ZrQtGQlUUm3gk5jMDlnllAOPfwm09mPo1iz4UV4thEf0LuxPPApvqy1Jsvv95tug
CMkoZfeF9uc7O/VnXdJkoUoS/yPZKv2yZQcjDMsW/opvLQnzsHWhaOY7TS8W60ge
jb3A++gzLcbzGQkbPGBB9Is0gY7zW+r+GSIGOZfKnEEgW1vKhJucLk/14xq9ueNm
Ry91wlAGxShbjIHjCgbt1nqgrWw6Zauz7e3Yjw6Y0nToBOrAzxtkvd6E0572SX6j
fKSHbwxMFxiTOAz6iTVYYncsJlAXQ8INmnZcGiRTFrntRj91R9krzFgHiJfc0EP7
gzdmithRZV81r82Z4efx01DKDvZJAaKmyVYcPWAf0/sfKOxE0Uu9lSj9NnVw7r5n
WUe09msR2sYcakmWFjnPBXRV0NDyI7IuxAl8g747ksA9MSCmgJILt90uJFv3Yuj+
j0+M3EUFVSSp1RMkrviGpeOZK+5XSVLPIMB5Ple7FbbXhuzEHfiRoJlQDwqSxS2s
Gxs16pis3TizMmYQxvAMeW+lirenPVnt0cyb24nCcgsUJ/U41QSkQlB7C5TjD0lm
o1wGeBh7PNataVjKKK5lgnC2gYNTv0Sybxn1qWgp+R2d54aX9SrMfOJxnUKdqFLq
QYQ51Le1bve85UWnZePzoIzMGb7zznnbaTbn18pRwGGKr9YMXMQfhY9QS/jgS+to
6oVn9B/1RDNBpm2PWVPsOGl60HvfU1P8spncneu+zkCpsbC6eHHTQD8nCLMxxRDn
4rBfT/09JF80hhi8vGhkQw4k3QEhApiIu+IK91WU61v5SgCG9ncHsFtI5L/ZEocX
eHKVHx9Z4tkHwhcQJ7iHz6ElPP2aHt5kSrB5MxBZFyoxY4SyKdGXv9adVQGNNeOn
uJHFuqcD2P0qjK1davdSwTI6S1d7T6MyIltymy5Uhfxnc3IAb3VQY0iQm8GmNAvd
PVMC6DM0bU0wx1eNBi1KWnpK9M2UQHRByQ+MJDKeJpC1PMODmUPSXUo6Yb2V3qkp
amYmBALr+wVpQjZ+kQKhkQCrT4Ma+DlrkstmaLMdLN5Re5IFHScrnfT9T2F2hyvx
zssJLFkJBfbjk0hQUFGSizoYI4T+MHxaetcVJK26KYxELIGDd1vqpWufftEM4XLn
8UFYIKXf1EbM69UNlaLwGZ2J6HywK+oeApgMgd4HixfurD/oeeHBXfX+qCsNEMSc
eHYzLhQOFBb5cz5ZY6xRL1zi+z683ItkE42FT5NZRzSk9KE9BysvqPXOBK41Jz37
x9N2Ewxbgyv3eJMrNsipfW4qWgsRztqkLSBVz1uGw2dI4t8Slc3mujBydgnc9gAC
PS0TxPdj5Iq8dhwC2TR6mf2KNqQeb4N1HvcPYrbpDS/IxlC8C7YYRELC1qIO8j9j
pLtTTU/M6Aikwa+eY1f50OfUN2S9B4QoooXul00h9fLBjfz6o8AghFZPPLkRxS5J
QNtHNGjnfv75y6hrMdl6eSSMx+rwjltnJBVlU2OtVF1pCetNJ8pQtBl6ROkvvv4l
DpIDQqbigBKghnyac9VhBSQjn8eVN7dBFR4LC/eI2ttwO02c7yhwFBkHjBRIgcbN
31qOYhHH8mmqM/1h4WWbSrSj1e93GYtAd53x5Ng0YIRYO8HJQIeibiBmGuxgeiYE
cZ17IY2GNOOliIStm/tLn8Dct40v7sPdUdtfuWcPKuniI6MFnmTyIYGaMqTaMtqz
uxplyyhGscBYKGX9RpNZettM5zvzD+QewceVjrb0C5Cdjv/Sjv7vmJJVHi4oUEIO
FMcl8R+yaDJ8zcoIoiGFGdhpWlYEEnUlJll5FgQ2gvgOVCHICBfrBceBXT92zhmq
udVk3nq4aaiJa79ZAvCG0Ckz1NOM8CrEuBt1mWmjDHmQIgybbOG1OeUawabrzJHl
eEe+G3ggY1W+IEGSaCPPVOB+1jEPs00s5C+mOMWfSBaqSXuqqkOvSZlnzm0WCyIG
4EUgqhrjtQEaLpu5KUPbYoRnNFFOVbmIbX3eSe17CdkF1tXVY4Q939/KMmAIeqdl
hD/44Zzq9WhTX0TGrL2qCyRHhYCRcR6qRFWm3bGgdWI6a9+BbpXQZdrjd9ALVQ3Z
bp2dsuXjOPbxbO9X1Ld8oPwPAgMjjEyvzIynEPlCCSS21+dhnHXDAyy9JiAXYif2
0IYxjohbeoCbZAtjd7SBO7y3nz6dRA5naynLbvODD7vnbqizN6ipicGUyDdjQ/9Q
xeH8Jktk/RWMeEclf5Rn5ttFk/qSNTSRRMoRSIiQwsJzea59KlVEmegnPP6kVGQM
2tM6ntlfiiJiE7REFX9cgdKWclPWN4g+sTd80t4UNzRs7WcnHXv40/JuE3NnNHTv
2Jgn5Ll/rtRln9qbWT+kcKsNYRBeKVx77zm8UsfqtRUDE6qLM0gHbO5ZUGYgA40A
kvBfIvsQRo56lnkyfIfaT1ba0R9y+NPmQaEwo8xobcrvNvO23JUM+OFVEAUGMjPa
zGHyTR0ccxhlwXjtNXKRL4D142UYPNbaZOZWGsUl7cowp3kIJMJz1WajNLFCvpxR
NYgEghvYrLMY9U+mGgbAjbZ+m5c10zjxZfZbGNjYFw7cI3prp/ET+BX3WZSp2uNX
+5JnxK5ADzLEmLyXzyExWfaDIewGJLd7b2m23di7In6HQ/YvW33GlQ48lu6spYyt
vG1Mu4vfjEwfYyJL9a7BxMPwo+IFe5vaVY2KswrQHJGP9MtrX/dwLdTdzK4srF+Y
OfeK+AzqMd2kC5QqK9i5FBbmZpgvP/R1chZ7QbMXutwOrYzt12Hur7EYZxPnDe/9
guSZfNOsdMSUL7jV5Cd0QkfrJePijhRAlhnClURLxreA2pAhtaR7REGZV37fH3qn
jRVWxqiT0il3w0MY9CCbo2UTyDJHpeGnG1O7EnH2xMWSuf1pCmjPZKcPA+6LMJyC
HzZjHirlFtnQW47Xaw2DeHsfWZ9Uz1YAUonXVJMhisjlsZnYnvuxDgygkpR08wuc
xRSmGtuQe4PuV5gonfn4PrUbKSWL7XxLaiAN3fK8r9OXyD7iy8vVOkbvrDUaExMG
7XUMbY769MEYtOZiQ7RJkbeelsdbQWPs6dV8bb9vyFZXGUtrrkjhDwr0x+KrXCD9
ZNYLh4UdypIcu8YcXpWtaeC1zPLETxhH9Y2Lz4hyhMcx8dj7+7Ih9/wxC0R8RmKr
NQL2JWAYDeU0z9LfizeqJhVDyFOmxIioVgN68GwewDGzmZbZacXyFe3xfQ3teSg2
yAhdd7xo8aKu89SafIj5c9SSBcDH8tMtYOkOxyTMTq7Feba6KJtVwjPD8IB3FudP
OSob4YUGy9j6T8nR03iKyu/GVbxVWoBzV8IFrQFPn1jyEk7G7Eo3N+En9EGZNh0k
Zuf0vs3wsX/kTm+iTYn+MG+IkvBfFulznI3OEj8UzH0TNzKhV9YimadnbqLTyOsb
IGU3TyvagmWlwY1rS2mfpvWRC1/KVqQrlLXS3WnYVeX4nO+Lzb/itucJvzf/mohq
BlxNFDqN6tDSDotaIGfKmJzbSKfhV9daFQEYoBaOmT3ERdzV9RcYIhDRtW9VBbXm
L57i3EsXBJ2P0QRvaQGpZWrGWKSHCUdXEse3C1a6+jqWK9oY+UYvWSLB+GqrMe+H
HK+KZkPsbHnICzguLPOIA8Ui7K0eLRGBVxAgRzYeXQr/b4S8iEpupT8nC3+vHI6l
NS2o++Vs/aR69cXvDm9HyABJqrAt45pQNfMTg6lSn5qW+pHB2bLtaRxJgZjx1+r6
qH6P2IbvltVJLehF/x1b2AhC0dRfaKuEYDBwf+LvQnO/ItIB0+iLa529/1t7r0qu
ZuH7ZhXSJ6//obfApOUy+zMBOsIAMOQTDqPWM4q7zMtkqSpGB17e7YMRrA9yqJpL
BQinGWPEhAItTE1huwOOkFiNoSrnPMzuC3HZSBSe3yKCYCWk5PdW9eo9xTITz8wi
snDRRL4PRRcj9KWyu4hr0HtarhswvnyFH6Xxm9fh+glE1E7cBw1nLkBMcX7Uh0OJ
qb/HHZilSok8GF7FSOqD9eNXEu+VxNIxySFraaIOywaQY2L3z/6YY/pYMRQKtiLL
44UxodGHkkBBwITXT5qsS3sBGTfICYXNgw2Zocc2t+pSaLQhFXDUpOHrhHR8FZSq
la7rvOp7yoOypnUuQopXv1pz5uPuEAWwMEYx5v/6fwBXbJsbYXBXYTRlc5YhYXYz
rCSQ/kyYetFTim7mlT2360/WRJmGou9xnxSdmqh+8wDTyuuaJgDA7PghflWUsMW2
Ac9rmmaUXMIQhdXcOD3QR/ZVjaEdBc9gXqjqxqAQPYdhMhyZCE6btvxp8HtUske3
r4WYacRdDoSfHFWIZSLJsvSXUzv1YbfPJhtbiyfIIxWFlH0hu3eSJdCOBdJd4XEs
BSQTnLWvCTzbY3+I68gPnox0/ivstHggsCtvp4qZjIsJkBuKefKSNp2X+I2rbmCx
+B5uPCQeacLjUAGuVjycYcd9C6DUr7I6LlzTB70l/QR2OZeYoNXIxOtzx8cRXE65
1y9OQJQ69bomQFV2WVileqqbWt4XGSyt2o/lMkjqVbsVY8dOM487F7Z0CD06j4Vl
2vMjfZo7vYnu6EoepyrXo07XznD+2XB/ILxoyCeoFIjQCMoA6WLm6WD87tdHhzgz
HI7GqJa8BbkL8ah6Xg7AWz24t8A5lGu6wOgGh3Oz0EiBqO0+2TVxjcNdUdkswmvm
XOFl2+z6GJd/oQPFuvXVESpxRr99jzdd4GdOE+GyH8MfZMi1MH3lUczssiXQnqw5
nBvLZY77GVxK3y03YU6KYb2ewUacnKjw2TSoKykzCHzuPvSw2/8MZHfhTL1aa+Xz
uQek0+j9mj8C+yJdgj3w47nMqnHEwwPXjDa+SOzcjOB9M6z19iN/+UhYIzqAq8h2
cEAe/5VZuOW2Idkr+R/F44VR6Vo/lRjYFEgvEjjqa3xYVT+Q+cggxTtcx52/jB/E
L8Hpa7gKRSXXAH78xZ+7yjwwL7G9FYhZc7xQIsp2awI8yDRsIa98uaJvsZlk7apq
L3qBWsz5lwlMRM+TvJ417VHIQd3WTxERg5hod2obXwwlMLIfiFJXms50dk/6AXo6
9lbXH6fAt9xFJtRBGkHlUncc/ELG5V2iIR1E7QQeSJiFbaj75Ha4NSp2q5crkMcP
EONX3Wv+xEJwOOanZGrxLqZbqpvmVfXS5UEvwRX43nEsCGNEA0iJU/gQTQ/0HIvL
qseUtcAAy/piLLhqQvWdNhabXcgnieRCGl38/Dvh8nUN+Xf0OI00odssjvtWb2nI
NPnaVTMutLyg0BkJfYekj/LH+GmM47jh5nmmKDdHu/czxmRXRPzEuyWV2iHgvBuS
vnhlk5TviHUrZMcYVu05/Me/cWivQ/Y581eaTsRFk1+ZQ4zTxC1rI+6+H1daQ5lQ
rae8u+LqLsTX+dxjaGcqXr4ykHDNQMUy7xLSO/v7tS3aVwmnEiCZNHe+kyPc8vKn
d1s+6bh7cZymoDcYNG5ueBzDQmiwXBFFqj/AjVjXh1hkHfmtUpbGDNF0GuSpqR/5
uWvQ+p8mIgiZW401NDaMKXqM+hmYD1qMy9Xrsdk6AnxjLd2A6A+FwpCOBfEr42lv
LqWM+AR8UwPkKNTqGD8B4R36VKXp+9bXB/KjxYiXelTDk7bh7d/CKQmzeIlHwJh1
sX8+KRJdWcplyGhYFFjiTKqFVPghpJZ6kHlmGiq5auhIMYEnHZ9YCXymUOX/f6zw
5tXpR6bJzju20onGtblINeyX2Lo5hXBGbfLqX+YhTqOX7rdoepNiawxpPDy/zSAe
s8FyVrsmFbWOiMwUb+P6Ob9lRWtdE/wJaS+kYJUSsqyb9YVFFd3je8A2CjW9wChF
6SPVzasla7jd370KjUzT61ha/D8taOYho0vDIkjyNHRi9fz4o9Kb/yIxujpdBY0+
oF2AVI+MyfTdkIKrbv4ll8Yzj98Fp8BWOVir4vwGEnV+U8g3P6bPLkZEOmJ57LBK
WSOaE7tADvxCe7vVjykzeDqwRj4ph507IoAFSG6gWwmBtzhX4GH5uxDoQdyD+d27
7sqF7Qhb4EDOYznu+VTSGLqHiykW9TY6e45SYI8oFhOgkb94oFzClBkV+VNeRScu
CMK09rzHPCLn4ysmajVT1rfZYVYhUW4IVx45LYtspvdynmqksdZLyS12alAGdYiG
clrxja9GX8yCd9AQZ/uELmtSYtTOjkPqxmjLN4Ml4g3rD5MPI4Jcs/4+giPiDnUm
+jvIR5JaKjn1cmhB2YC1ArezKDhuzSBSBsgFaaouvJLC8qmNDcbPyrZ3zs/161/v
fE90jYCRICvk8pJtNmL/kKDJGG7llRBAWSRunPZWu6P3s+BhfKLSozbYCsEkBMTZ
NlJ5d6+huj56N9g0g6AWRMkd6UXaOA95f2VJJ0uCQUdB0zk0n+wjVyxzwMe/lmYj
7yIHg/NPZffKKIv95RWT6qYJEnDH0CPbKMIe77RN/avOIQ9sQOTnMv8ImOtsvA8F
ISOZskKz5LJEnW4w7F6MWmqqheGzp3IIMvqBVKtdSpxHtEquhL2hngr12JOWkNPC
PnbAtTZiZZ0tQP/xonElslEuK1EZoqDIE+tGpo4IlhtYSpyy/ul5ZHFA0oTDkdSO
d6Z8ihTlR//de9POMzF5SEZw3BaQZmTQ8TV+WfYZFLSCnLqeZFAJ5hXMzMBvjoM+
usxrr5pvF9DYXyPshqwVIJqa99Ydv0zsPpLtl+LVFlDfoSttjVSYQiUYrpI7I5WW
R4LrtIFa5cuqrZoYg/WEN9GejVWNmtVD9llc9kG/+rUBZm2gfyjM6l67b0gbCJKP
FpwBn3iGw2Seu69tDX4nC9P2ukFTV+e4gdfaogU8XvKD2mnXJ+1S6yHAsKSiygk9
vfLzDn6Vb/I+bBtEHHtm9uls3tHnLtCtqDKLJ2CYD8HOTD1upXgXL4mByMnX8wfa
HYw03/66+A/K6AG+AuG/c1wwId8G+VxM7kvu/u9OTeGnBGpJXtk4p+CJXj388umK
ASrsJ4mpYs+IBIDoG6kuvdfshpftvEQw6TQD1N6ar0PzmN+ZzivN/T4EOcKhai9k
8NCL9goIsolbrgWSyOXOuapM+U4Tuke14gPfFTyHtl1FZvIb/zFkCuTnCdbGe/so
148q5dLfbwOM1jq23mx46jJq/+hwvetGCrRpHTV+2RxYRWLSCswVuQMlK/mnpI8e
ldLgK++jcdQ90tqqb+J2rjr80CfrQ++SnPtLkvlhECdQmrVjx3PBnuwm4u4jAx9S
xEx1BIf5fJS/dF3BClj8XS/kQjkPWWOGQzYNID6xbhO98oyJ7ImNQGoKuMIGCSx0
Zy3S/GgrHzRwonPyfzj7OGNztv/YW8SO0hRE/6ICFwuf7HwFcQrP0erl8s8yCIVu
+GgTC+etQVx/MMysm7weXpdMOE312oJvIXsBYrdqYsNNQd5ME7lWUUEP65Tu1yLY
APDJRt+tt2ANqd+4+0+du74ezCXHEmHltMbg8sll2WOi2xUZzUC6qs2GoGxvzuCD
xarcWG8GAivot//D3lnIsp4xXPWrWE783URu06eP4FSKkoScQ5Y5YjkLExOTGhCb
fgNCpXu6TDNSrQTEBId407IHG5kueNYBtpRlgTCr1ZuYrXpGYYDaml6Yktk45x4U
4AJ2wVXZfSYHCGpDDAccgzlMZJGId+61DV6vJg+S2FMSxyHqU5umjAtfUEi1DGn6
2aBAWMyNKNT69vB/Gyf1kZeljLVlozFPINv8LAnPTaQpfZU5K8pe27my13M+UE9y
oKJb8yIctbV4pE9rC9gigm/Ql3sLibRNyUPW90eO4TqOmbMyatdYNICP5Y7obC39
bds22dNlOmVoYnGlOP/Ih4H5v+h1wu77nRT9eeEaZK+lpRbEQI+GETiKg0Vg8EbF
M7lGKlqZH+8dKNxo1zgFH0NjioVT8ZStoMYX4WGEn6iZPww4fe6iO2/EhXBFTyWG
QVgArF1/PyxdUol6d+ioMclKb4cbX6jdArqUWxnbm+lFVwW5myzCtw0jP3IHIOn5
Hwfbp10tDyfvabOrZhB+reDknSRmB2omQP+fJl55g5SRonksqWhCCXjLfawQwD3E
bFH60WED8Myjl8gtpBC8xncGeoQG5XdbdJx9ZuqHqVboB4oj8etTvPPrsKc4tEoS
vRu4tPPrapY1X0job3dD5YXh3MK8wJnyWi69c0Zzt37SwcRKmUWSEfqwyT2n5uz+
yrRFoCvnb1DdsoqqLhEtDF4FMFTzj0h4U/k21/e+Y8XgOv+IVeJWCJN8fwAfe1+n
v5zn/t8DKE1UZuQ9s//KZKTr+ImgKLG+brf/9ZL3HJp2uiWy+r+H2JvgWtgY9pPp
fOzumBcRYMaC+UZg+bBi58P6UEPxZNHjXYukPciqCTfXPzJaE5GA1plN3EMM4KDx
Kt1cZ5RyeWoHLnxEVd8TC3iUW068AaUII08V4IgCKiNTjcQ3/0y0QuaJ9e/dhyuB
DLJ+qSvkz6K8luUBJ/hwbTYhhTph4hJhe/OCbo7KV3tnSs3+HykWgQ3LE0CHjyVv
5cHXBqehZBdSozBsJLjSdQRlZo7D3eBtNdx4nipUFbxmwVbPmZ6sakvmVDPNaxv4
8TadhrCmAQVmAQ8FeOsYuvhZhp0/Z2cuhSWXwp3GbF5Aeq6fFLdoGNDhnuVymVhC
blETU7Oq8R6MX7cUKgAITTOfrw9+G+XnL4QgNE3vmByxlHlji9Xk8FhO3rESBr9R
8dNJhfsi4gzjU2gMsUkNXNQ00WFMA+8UL5BF9MIfSBZnmviWUmZpTp0YzdgLx5v1
Een03EHPlVEwbGqc4hojHpJVJz0SXzI2oynGNPk3sSqyLEjklR1HVyubD7O6V2FX
RrnLsIeSGb74fGki6nnxx8jOzfAB4QGQ6ulu6DbjCX4dbx6vDjJ6jihE0sSi8hf4
m1SJ2B9d4GacwRR7B7S2yaKkhIPcjWbbAFeoso/terh63x6VdWF7e1twuSTeS5NG
ygq+IatC0wLGNjjQXTjSxNbmSDvYs/Vz4Gzwh5J9nvLyFjJ+jvzHAiUZlcLZDBrv
rB51naSnEU9uznS6hXUqyb6w2JvARUUK9mqP/W4CnnsU4X5RXqXAjAikcJbXDAvc
WNG9i9bh7fM6BNXeP/WVRo8O8tZOFaeRUy6D7Qzr6qX5Ia5zCaiKDskSBAo2W24Z
ui9WuTlxcuOZmdvOknQLgoU3N3bpGU8XBj9dNEcmPuIFN14GS5I2rlw3M9X9zYAw
r6kJ/RFtk//Yz46lcBMz4AQItmRRQUUvDZgxFCKQG2fEf1/5u2zAWBSKeFMHejO6
AwHKI0ek8Co6h2zIYS+a3iWeyFFVjYmFEghvlqI/fd7N8I+AVB2zi+BvP3eC/Q8Z
JlRidcfZ3bEkgWFdz6phbp09GEEjpyPEQQ0KcDkw7io9YNyioHIRqySGqo0XiwHh
UqmFjVEbu7uQXSMqhcoPGqcPc4HU6NJFFPS4aAuL2VIa3crIAoaJg3LIaW79QOqG
bDjHvI/l9QOa1ddUwjpsRPkfR06Mw+WwBpsngJFBrjHw6mh92+mQXEZHmMQ+BpDB
LlsF6yUJNd+iSiM5/VDNUBWSyatxvJXR8mRGRDv3dRpX7DjkzIAB5XJGg0v0Get+
AW02Srcsnb9iJSZn5ENfNkw2z+bCBe257UmaH3f60m/vbOiVD+8koktGmtg6QQVD
OetPjFg9K2VUBH4dVemX2/MaD6kRei4XU5f6Z8W9YCzwAaroE11TdEMaLoacqxHv
9TDtLkjFedofiZhli4bLBrqCDOLVQfwtXTnsplqhjpjNLHmG3GNIrb+QfSfSt/aA
FlQo0fc3X9uOuyoYYBiUz8H7dBonZQjK2ghAQI4izUQs1JA6+ZT3hcbMiSwbBjq0
K6Rt3T8Us6d2KZYL0kCIfPnkF7SgUYS0W73oUP5IVMK5n7SqrC2R2/E3omewN82Z
JgUBns/cKEgDIotk9w5pyLgnCEXw5cguiFcXLm0TeqXYmqHtb1wMb43WapOIlnmx
E29YgeIGxKw5HVfINx4zJZmh2zo0De+ZqUewaCaGWQTNhWXaKA0gBD04Yi0U2+ws
5uEHmg91DydOSi/D2CQA4gJs5Pnmg9LQT3P35FJzpj8I3kPM/k4hD+DHjXT8cUM2
nsUR9eF7VEbiQRwBXcOxlhFcm5DirTqAsdnphIUCstVWymm/0m/JliVL0DUloPS8
8aK3yzYl6wd6xOLPIaPXq5f+rggOLAuNKXG9JIdnTLuAhEzC1cTJPyy5a8ip9H23
gRtT+g5xCPyumd4NsBz9bK1yJqznI5wtBExW9/G5AZuBAOTK/bem56FRpgYf5SYP
X+NANgioSnBxTqHyIHce9P9S7uYIf9xH8o+KcU2UEn3pFDct/zK0+vQs5B1YJb5O
wRSwvBR4du6qK9SV/Co512WZpEllZirng/6Fapm6hyOhLedmuB5D9KI47UEk5hIO
28ud/MxKmMM5CU9bj0QmgOoQ6DPq/g1QmmlB51FCwG4B7I2R2d5CNmkCKzF96/8s
AvND6JVKqVPwmpJ4J3mkNXQFZ6SFmUVSM+XG3YOkTHZv4Wx9+6Uluv2GV0tWwgvs
SDxrBp/MBK/7LgYw0AwW79t+31N3sM48u6T2b2qKl8cbkUcJXLTsV26J2gHZj75F
eKTgH9yu3F8BwKgyjcLSEVHaS5KNjNV/CUX1qwDB3fQKyOH4VWgB4rDqto6U5Ao8
UYWRDy3EoTOQH9/lTWYI9lY+gE0V1SpWPph3vTIksk9wSosSCl7TMROqlGKjlGLg
8cd9xZeWo6OQlh91hKaPLJZH3JYyPzYZpQjkKN8WjwoHKh/sE5VlQLBIDUG3CTDC
W3AJZ7Pzpc2MB3ba23i6L5RRDK7egmR83RfAKu4OH5lYTotrv53VavH1wauPacF8
q01Oor5KCMNW88LPq3eaSEzZyVlqPCmM3XBDYeocYHE+t09fhJOJor9665Kclz3E
+WXlTWs4/LGCb1Pq/EpR39D9BwD7paRGfdAO2dKX53EN2QP95z+NEYcSh500M1V7
Ust2ZAwNGByQuAiAh1PFb+Sj12ywt18uhX7Swx1QKMUfTFpAOEXICCbFO/cnzZ3V
+uPKgks7kfvH6Wn52kaikwbDgJBQEehtBJBdzt7/9GaUJOt/KH1MaYXGbaxQ+9eA
EC9N8z3RZR6mrFEDe6fpKwzco2b7+iwaT5bvwHHyYKIV8IA0IH2406m74GnpOr6c
njIQcR7kmNkB4y473k7d3HBXyLkYupV4zhEYvCXB4u3TLEUdNe3JZZ+SrZfE3pPl
Ezflk3oUHL33Fc77nkvaSucQprHSTYJZ3s28dndA4aMTWDrlyJA9wzON+oE0TcVw
xAbqglfaI83GFvdK3XAphgb3ZDv3EtHftmevMqg/RjPvf8feVy6PgbwUt3WbHXfe
WsuctonR4MkN8YCjnFcDbcU8N2BdcjwVxfTDTNMZZPZmhcOIXpPeAJcdV/MAWc+k
YFLbnPwzbs0cKG0MD3LFY5SapNsf1eI1kZF2NREgsB1xVHtXLaFKcKrYvXyCcXjm
fAU1UiSC8L+CVGLk8CFmiUa1MeZWSk1jRcSaDSiNOSe1/PgLGku1/BEtePSoa7W0
iy/Xj7w6yHtFA6n43NvdT0Q1pUwHeaWBH57mOMOl4kJ8i5TEsVQ6vj0ZXLHHIEuf
0MMS5Du7UuhbMxCbTPtVxQoQzV59MF++eJ2g5PdTu1edOQ9kOB7J6ntUavTbLgxb
WNlV2hxMZXVvIRPBAI1kGvCfVCulq31z34UkTex2PkLH+l9Pk2P+WNndU/F4SseA
VnyKHqSueZsXHvDil9lIKO1ZamzbXW1j29u1rqQ5j4iqY3PuR+VaMvJcb4ewb38M
bj9IDibYSMdU5ZANvuZFLr1QphjSGNX2StDI4jZ2oCIttZeyBUvSDujB1NSpTb41
6XmqHH1P2kt5vEMBYGc/nUhHUqY6oWmGbh43+yeepSFGMRZvvFUJMVpgXrqIQlRH
COqKPqrQh+2PXx/nkaBUMHQM9gXQEFW2rJwKzDyCHMK+68gJgev6L4VuSzETrkVO
hGhHhdyDWcWkh8QabjZY41StF47u8+GKe7TqIT8SQQfMr50zF5xq353HitekbtSB
Mb7z2UXh0vQst7ohPfwRreo5kvAgdT+W6rOY8ClWAezmuUG9+cToVC+qZb3yeynO
JMvsrsIOFKtGELsS7OZrkVMUJU6DqNQj6Eo18MDAeBh4f9cd35L2pCFuJXLxPrS9
p++aMeodIGm3EOc23wZwXj+tBLtN04KEQjgo1avVbSypfoLI/xbz6piWFiUiyXXK
CT1dchP9GXDSrt5i/EnF0FNklfS0C85GH9tAt5qOsYj415wwC0r3vNMLinSwqdxI
BJ69BxWdq9Trz07CkSAhba6njXDSn9bJsyZV/GF+VI8RM/3RdssEkx//ZT51Ji5H
mNx+QnWVCk4vSbmtt/1eOI8mVr21w/W1AFqKF+tKz7oQj/ntBiqC4skoM7Ojn61H
MyK725R6wqFdjxhBOz9tCRBjZW7AN5UvymBrPJjkV1f7HxpCvrwS7GpyrfxjYlAa
GECXskqKnClVI80XB3ofcC05AvuI25ybgngTmQ1VBsfP8jiXdc5sP0yWaf0XTGCW
O7IrwSamrTReIFu2O/BLmN63/JnD9DEGA8S3uUrGHJMrSRQSMd2iMBGe0I2cRIVc
hips344EwJAlGfCgye+N35xNqFBn3rQ6fxjD+RtDZYxC53JFO7Z7UzKty4O8g8qB
RUlZDne/WegNIW6YGKek5ZWU0c7M0vO74rhWhS91Ch9I63E/MWhtcrso+0qjo8RT
pxHy6s3TR9iAZVCgb45vjmmJgPaV2PqnMDrz9rmxpFPDdJKaOqQAr6XdWxY22Ago
WLz3MegWNluj1jxPmF9M2wOTdkcSevEzAg4i6m4phx2Q/hm3ZzAWxkLuwScURhN5
O9347ECmMv8wVBFCTAwnc9DHIw2LgR7asAaQnwKc3538SCvLbTPsu0dUNQtbFtZR
2stlYk3V6+MYyjGpJo45nBVLRAcFZ7rvZ2RQnpbWykohelXBb+L5kU9ghluObyvd
1oTVF5b5FCw7n1sy3aqtDMxCY7+OInsPaPCP5BU9oeurj0IfSHdLQXB1Xwe7JhyE
OZyVASXFK3n71IxmRWlgVCwWl4TNudNteNkTP+3M8LV4ucnyOFZwsLQ2XzKngGa3
RyfRQWpjP9Xofhg7xCYr0/MLmPEo/E2Izk/wN1n58gAy/81GZresy1UBUXsU/RwQ
saUZ6ozMv60VvO/WWrgAIzQkGCvSAhsunuIUMTpf12QxTgAkccTJpFvuOj8daSSU
pq8gE5U7cJNTKSHpn76fMbTXzxZcyR2QUbiuy0COzeU0f/F5XkkD1vVe6ULO54jn
kTWRfZcJGHYoAqoqJ9AOExDXz4sm+DgKUDcEOhW/wovzslcSiFJ9cufcIMTm6sFh
wBv3Pq2e944lm2dMwZHWbG8mHIbroWJvNVuvILXZYrnESNiu7sVUyFsGATMrMOWb
ZYMUZKHU77Qd/72XUIF83Qm9ZiLZBwL+0jnOskUQE0bkBzUY/4WreqYFZ/iKCvsC
bVJmeCmX9G023izc6W+/wv9AMH33tjQ3XdCgeWqsfICAVCfYAoKJ6/tT/dd5yEUH
6fd5FrutjQfJGOKD4pc1mdT6DPf0S0BgsDu2OUa+3XUR8BT6kpgVtDvpdh4f+EKC
ZkPSt66trcf698wF6Krwxe5NY6QUDnCHTfRSPIRECYbmwG9uCs62h6Q/pFIXwhxW
dHSrL0xPItxjpb2aAqWvtJEuYViR79HSXnvUnKRkeJffGtxnwsySnb6NLUf8sv7g
C8YPE1U9GruSxjr79f7GRD8FTEMozZQQzpFiy/uagCD8ThM0Sve9Qejn1MBKXyjb
90je0OSNeKhdLk56not68JlWV3opAKlvNz5L4zHf0hmmXNwzk61+tTEw4jh+1Jm5
K1ajwa7apvknXG9V6JixhBkKRWKgnAE0okzf9jKXo7Wj3vUSTQfCmuZdDms2y0LG
Xro6qtGpjaxxY14RuUsUt7rVmn8ir5HIjA8RhjwL9eacfR6G2Hlc7CXBow5m1y3W
i+YP4lXXAg29SuNieOxdzxtcWXa8EDBZeDfvEgLzsQSQXBtF9yRijrsgT9fHujnZ
UdFlTwcHGIW5zdODjlw0yRKCOa0vVK0wM7RA4XOACaHM6PmrzYmLRBZSQvOOUdar
us2LkZJb7LLrzAmj8N0dVJtQ13zxQGk/LydIeE8bXm0GwCXhCJHlwCd+o/vhWU4B
EKNEvHBrAdt9YT0N1uqrjtipbZ2neDDVfZYyspM+4Qo+P2ohv0oKh3k7/BkK9tK4
QcSDara0B+mutGt+J/BiMqhJKGwKUmbsYUnHmuYPQpd/xKsEW2CSb4FTIEKqpEjC
sG9ovO25TZvhuNehc1wecF4YLdf94HZCTW9xiwcadm1/405yMg4B5VIw4FfqHX16
7paDkQZRw+OT8CeWcia5DK2+OGLW6nAoWblh+V/RY/wK4T3g2Wcmwtdo+cKKQKG3
fFv5pfjdKk0FXigKJ97kkRS0ZLycnDsb89pBgt+PhbKDKYpUnnEFKqD5CtXnOFxm
pnsxoNIlX3n9zsTzobHXsOPGMfoeF61OlSBTwIlXR1lGWPe8P7mWXVi7tYq7XHDU
5YfS4MWVGCnSFr8xkMK3gYpTEgyu4CpkiWnBzbj/BMRx+8M/8Cbux5DtuF+G8WMd
KUVnXIGQjNWecOj7B2XeXAcV+BJkYyWKrtbZwBdQ1c2kuQIeoLnfB0QBkGiBUlFy
C94C7d8mR0ic/aINdbPN/W5ySeNH5KZ0kvOrcyLU6sa24LMRtkiYcvbl7u6sXAuX
WwK8+2X5NxFKENKAl8N3zA72asCC2W7sAPxB+hoETnvvmmxYmgEJ3T+B8AyZ7NVr
/4jhcMLmhslmSt0ENOVoAAfXsMBSQSb1jx+2+TR4JsWbL1NYSmmQ8Skca1RCIeSQ
6v03EpGxviBZnj6gg8rdqxoTjrxD8s6BWffpZR6QU3b2pMM9yxXPRjsaN+Y8MShB
tzAX12uRckgxAB5E7aVoIBwvO9r30LLKEKx+1TAUeySQ0u5kduOTI4yjPl5ZxIX5
tCBAF/rg/ZVJVs+5y7yTNadDr4paLqWbzCQ4Eb/0DBG18GNknf/bNA46I1NukrSJ
+f/UNln9fq2Y4Ye/YKeDv2yyZrDd7rpTr2dH7oS2svUsdlaCsTSWimCqp/+V5kCu
3QxWXCQCxWHnlg8j3Y1pWY/kwZMgPB2zHk+D1KgE3M2QLXXuu12iC9IpI/KIdDwc
ebYKqCswU+aD0N1i6lMea6/ARig51QiF3Fk8CI72XYqvp9aVbnmohtLq+0qhXxgk
znmk+GCROwB0OabyUAWwXktGsaxdWPn999Oc436Ec9ObQCOhjWf14vMZI4rwN8Z9
hC4q1LUFLrhsMvRkN5F43TO6j3h+SejloKTwz/BT5Ycbd2TXEDBs4y0G2l2Kyu5n
K78SPDqFF1tBjA5KCnD6s8qA/QnMO4tfpFeGsrCpA4i6DTKfr2n9Xw0FTcZhtNlJ
Tq8E8B9xgKbKmKRFIvcjtRjyWMC+1x+cvG0EfwFNweAmLCYgXPUKTCxPW2puk/V2
rCvElh1Z9syOqai21Gah2V1CUPVRAgcnZZBBNzRxuENqVUmYrZ31WkgvjU6mzDrF
YYQopQCNzquSzm1CKxHWwEbla/FGbQvXT90F583kYvcTgF14WDwVsUrAiMq4Gg2f
svbXSL9depTR9EMTwJJL+lHE+2AGYMjdOTrywV4YSlIFR+KYQv/oahgRFgMwD2un
8ggLjPTIlK+YEEG97rInz0pvj1Uc6Vtnc6bW1T+cmIu4SU8dEznDUjalZal8w4x8
fX1ZS5hniq8mGPWrfF6CLE50khcnnn8l11bXxs3K9OL7pSLMcrbdJ//cVFZlySoI
m3oCaYCjPbGtg0YY8yAglxTwuZh40A8giaI80OFzLUwuhn6AUbCW77ZZ61WdjzbT
aEeQ0nNU4Pz4GRrcgmN0WC78Ko+wxh7O9G6KMwoc1PGah5vDkAj2uT4WXq3O1YhC
bgfMXcz/AJApgRDKXk1YBEer9BInQf7j1lgpSOA9uxRM3oAhKtQfjvgSBOYzbxbJ
AUyfQ27DoF5II5Vih7zDBG1qmIqgGXJmVTn21qTqvhq4BON7oMAB92bh//PNU8/q
IkHYvvwwQ81qYKTyxOunBgT4rNu1SqjjYNsyE9qWcEEteHKo82f89EVSEEzuHxf8
AKqdK9yEluDdOkXUFUEE91g6Dlv66vHFNeBlDOFHlOeUbN/K1bFWdJZm0+R6sST/
6SJW/nIuHnmJORK/iJP3G+GYsR1Y4UXhz/+i9hJD90qh7dDtlC4Vgfgd57Udh0f6
O4C9I3nRqGbmiiHm17n5j/7NiHGhwk4FvJdxMXV47BOJsTXT5/MCNjjIVXw12vPo
GXjy8xwaXwAuQsmxG7RX8/qElqblWjBN/bCZYWi7VvFJpoAp0z5be6jKlTm8Swlu
//pragma protect end_data_block
//pragma protect digest_block
PxKrmcqhMU4VakQYrwOf12u0kiU=
//pragma protect end_digest_block
//pragma protect end_protected
