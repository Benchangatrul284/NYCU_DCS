//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
HLKjwfuGM1swajpIeKRmjN9fR6Ieo5gkHEaXUxqG6qoMooOiRaZopxs21ompQLgO
iAy9GSr1Mp8AXUwOBJnMJgvlvmHZRt5VZHqwUVohbWcJWCqtfavBNVhB9nqndHac
WyeUQLEwHVBwm4j0qDf5hGwt7Fsc8GeDcko+zFIkwtbMffTCdXHAYQCJJoGDQXEV
3ZtHJg/ObDbtrV6UfbFRHAzmC2AGCcJWvHc5qBNhbAdAX7Dx16Wzl9ias0wXIuWC
TRtIK1SFzpoT9GnTcHn515HgcN+u10Ak3T2uGsPzH3j313oRADSUQPiAqn5BkcWg
bPHbl2jALdyQZfsDVtr1pg==
//pragma protect end_key_block
//pragma protect digest_block
WNM53dqvHD6CVEdYi10hi+98Am8=
//pragma protect end_digest_block
//pragma protect data_block
+TcOV/YP7tfGymfxmLF9LLvqBzAvNaiTklKORg2ny7TcNZCBlJCld1Bf7PqKM0l0
JmOaCtFgoNPW9NUvOIFBYg1yi641jPi+mQyYcGC2IsMHN6zKrmC0tgjrJneEaiCH
1syKZFCQ4k5qjq+eI4TTzuFhlc/z/ZHNcU9K5MOrpNOQOcnVSJMLhUuTQS5379Lk
W3d1rh/zSj8zdRrO4S0JVckYO2AP30BrwwPmHx6jMEaara/McP8OKFLQVRe9ZGZo
QFDln9JKdpxEplldN+WFv7ehk0W3ob8J1xFPatTKwSZeP6sysyxlyUOM0H8/ImKC
WnLmL0mmmErvyKR3kSX5gpCfMdB4+fJQK+GAcSLeYuYFO/1pAnf72msYsRw6msj8
OM5k1UOZ2I5sps3Wf0lAKEZcyNhdqeqrlP5pHL/SdhyCwlrK0xSW/vM1cxmpBdVK
JzMbQbqU5GWWQcaCEbfIOC6JoyZ9Q7tw/RQ2sQWs+XwCIBrzhmAhah5yjzJ5M9t1
AkwiIwFapu82Q5LC6PXLRjoQdDCZFrKaiyLHVM2m3jVKgxbbcJ8VFadQaeLoySV0
27LoXYvI/Pit8UN5Os3lUpuv5xjVjlCN/1yfzUyTDZ3hWZqu6rCKmu/BEFdL0OCC
lBI9nY/aiFIGwNrKbLKSVD4JdLmPUF8Nk2ZkdiMs0mlBZWfkHpKdqLeRriLHWrOU
tj92x+taIBpRCUEvBX8gp1HRQ2AEnHbcjqKJ8WrqpQC9gkaQulBFdd4ZmPle2q3v
a35Gnn55w0/D1IGRNDU7Omn5udVRZ/MHna+IXrBS1H+liKKac4Xf2xHumr2GZZSi
UyF6lAFH5yQfjj/Er2BSOk1i3Wnfr/pLSEkzzOF0AcYcj/xqp9aQoR1IlOi0OkKn
BlwbQMCirzx012la2NxuYH4Eo7PZNU06PnQ4Mf0LYNHO+nxfXY7El75TDCwScUwK
RIqm2mfCSk2oXHoPRfg0tb5Xj58wwWagi+JXKoYG9RbZNU+6U3872PIFyJb/wXfe
jMtzQ2GKiougzV+BADGnIhBIDeMHIvqANKmPbL9eOVYaffIEkWUk42ZnbYswpKea
PavifJPsEpLbnhjHN0GYZ2foTD2pYO/TmbEeSGr/Hv5bFYV8YJJZ9c4K0HZnxKCe
quOyXy7jC2aJTbFRw5y+XQWpxmcfvDJIf6C0HSS6frb6eLYebVOzkYxDPGmJ5PJN
LAeXrejVJABQJL8naox4VHXKBZltc5fTGogdnzvdA+iHwTpplZeYpYNdQzVKsq+v
onbd4U5mPhmilxl3tZuUHnyteN+DOP3xO4reYAcVhumNT9sHpvaD8m/M8kya5TW6
jbvMwbtaK2fV0G1KSvs28ZK4yZaQBawewF6J0nYAkN6hk0GZDYrhPr/1elXUYgtT
sFXYUKtaQu1EhDrqabwC9nWBCOapNO5UqpwjgXGQY9IRBnXakdtNw+VTm7nq+LxO
jqZI92vs2CWI4wf78A0dOfFApJUtmuncwChU8EXxdCUQkpczmycnOQIUIN3y5Odx
Z+j+owNi3uxCuLMtWoXnJRJ4FqOXJSwuv33l3hfyhvx5wLMdvJnyKoadM2mI4gWc
jJiP/THWu+SWoaYVCwe0ww0ijckOXryitY+L9F6RuOsZGyX7QFXLADP4K9N45hTJ
7pTjRr3X/WyZ0VD+HTVS81jPLRhWJksvJ/k/lvAaLJ3FYvHgVaGdwKp1wtbi4Gh1
FqItYQqGdRCN9urPPEHqTY690AiuoVQ7+pNERx01OMYTYLYhF9tpZLusj/uwiu0K
qiMroNNO6P1oUnYyuW5l59+VXLxGtpy93jyw4g2iwIe3i6KRIERHBooy4QagQiBQ
FwpMC20h8L8BzZ+1I43L8/QIFzESYu2NMY2GZlHQJYI=
//pragma protect end_data_block
//pragma protect digest_block
m4008U1TC7izq3n8Bl+N+IDUBvE=
//pragma protect end_digest_block
//pragma protect end_protected
