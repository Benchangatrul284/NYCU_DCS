`ifdef RTL
	`timescale 1ns/10ps
	`include "MIPS.sv"  
	`define CYCLE_TIME 3
`endif
`ifdef GATE
	`timescale 1ns/10ps
	`include "MIPS_SYN.v"
	`define CYCLE_TIME 3
`endif

//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
gkfcjK0gG/LgSqHt3eYniZ546ALIfOichcrbf1YHa7eGblwYMcpDB7sXJNfRrJz/
QkAm60Qrmd2HSra9bsHrFVkgiSCGzVYK4+JY1HHlbFGTXRSAdXQmbzwv9fGJAQ8f
gtZkysjSazeT9g9IjLq57LdNO1hMJyO0IKrKWNtheAaF77r3St7SCDI/6Ahhkw0G
dlFzNNS5wiRcB+1o36HFWGGUQT2ft1tto8iA14hWsb19WxYVO4wuzlhbA/ZPMor9
6WEHF3dQeLharKtjttc5GJeM3PdrL3VTjpDq/k9IIb66DL1pUq40cdXi4GNsEInC
Hqj4ExkuvagUHXP5EKh7Cw==
//pragma protect end_key_block
//pragma protect digest_block
mghiqu+jd8442xyFt0hMkecLzPY=
//pragma protect end_digest_block
//pragma protect data_block
EUXVJ034znskaJMNiMPzE5BHimmhdNrcfPjcOa0CN6C16BpKkCyrJCR79pJVH24E
4k9w/hFbQHQ5JcmfeFP4xrTXUNrFXYXbiDunq97Z5aBlXBzW+QfYcUvfYN2jqqPI
KWpOrpwKnnoGsGVn00pnlwEgpKYhehq3eC8/ZDvv7EI6kYxzyGft34n+Jn3F9BMc
UHW6lcf6xYdI15/DrhyAdvMror9ZkJ5HJ2JLSFm0Rbt9IvIFynavrqO54Rh6A9TL
hp/B0HhPYpIa+IICWMv19jWC0PPkqhCXaz7A12Q06mkd1P4VCOT/0/XPW8xqy4FI
mmcxPItN9Q1dy8XHdu23FkjB7xy0jhqZ3iUm3LGsRcPccEdVh6KRah/7Il2l2r6M
s9E+NO5t9KqeMOa9lNvdssDD3leVgAj/cr+rL+usrpsadxXw+GSSf0Rxu7Q16YJk
XYBdUiyE/zUtR1GcoRMyq7SzsIfTYvxVFSL/37gxpBwKjhqeCj+Dhx6nlkMbkwpj
vg7Np/EgZXKXQRKPmt3CKisyuzbJQsSFvXogBtO4Z31Upg0Ndk6GmWOMQT2oxFwn
rzG9JbbUOnK6A2N4y4P6qwcgFBUUyjapkNU1kKWDDpYh53lDCyo6ZA2f2almAuFp
pzYsu/hjRSz2mQLAjr/1KLyzhprRzMlNazCoyXBnG3NYsSR0AkktHgCeWqtzo/KB
scFDi2uviJjTuJfm8xWghnxsDdTJjplmYj2U3w0vrj49JPfY21foM4XeSvvsHk+j
VUTBx7IlzA0lwvByu8gMl1PBKqxyQWvSElckIqD7ufdgYiT74J+qjrsNlnjIkMPT
lJfQW2Cx2sbJLzpSCCOULjbtwOqaOXeL71lQSWaqjRpXzTd1oH3XZzk0jVB6oMUh
M6SY/MOhTxaM/D0mXXDiNY4DcJLJhokbiAfM4nLfovc4Q9GRNT9wpJnY7TQAcIl8
jj56ZRI7PY+7jWsvIoAbeuoctl0l1HuSdsZ1EZ0O+AG5p6dCxi4KupvAG/b+bD0E
gb4ylwregBA1uzTmHmXmnxnVnNzujODzriSWxymQ7hZE0quDuFn8KGL0ZKmhPQJp
/6mzrzhSfo5HjHYsai5kRqAZJT06S/W7QMm3q+8RdkqDuqqFbFCtTAtp7FI0ZShu
xHWt/zxBSh9irkKZGKGhRueKnL7B3aX/pWDpZjOQdVYSPGfT4cEp7eyVVFPalODU
bEdBvIpXF1hf98qYX57M4qR6/dfnRYwJ39mjxu1tbovsg8wfBoIxaAPMlbaanZYM
FBl7tf3tzly+U69kkdLFqB1yltueocJAIRolcId7L9Czv6govZCVyvCOXvvwOjn0
jgGfiNpn+9aokgctIQl8QCVD7MCQ3w1q1JJJ0Q7HGwgAsF8PtnJUoIioAhZVYBHw
jvQFbFrX1H/AmDEyDT406LEgTr0P9WzUUhR/DP1fiXX712Cn79AoXHTG29+FNLyu
YL1Txx5Hp6yIWd/tqra2m+Zd6laP74UafdVDFfs1HItqF0fibzLO29KhTzKKeRI2
Zu6wc114ZsHOLNQvS5swNSyj1PbUn6tSm67aXjsR3/F79fy8DCcb2+t0FcqyuiI1
NtgVYxfjZWhGyis0yCEEW5RpLrMsnA4U7HMKtto5NSN4TIibxlbXGqjxfE970q0q
WC/w5iOysZIPATcEOREAPnI/mbVhn8hLIvp2aj8ToVV4srX+1l/gdPbkyc/8zK+W
3Dg3tb/xv6AycWUP/TNGPFSvCCgnqOj0hZAeqUR6kIJeHPCpkrOR3VVpO8ZHpk8C
CwePcmrGPjRkcYiFqTYpVwkD2vEKtpRgnBK6cqt5d+qglznCA2wx1jt5+iCHXt8e
QzLcTUHog3JxEQmDlyN3g8fkxXtOxRPVunVV6JTkN++7A87XV/S3dC0GSclYyIyq
n96fow2akZvJSvt4zvMw2K3iX5FrA9ms7CAZvnISULJiAcTOr9mMG55alQQO+kVG
xicDP8weaAo+MIysXe9tKGXNNsFsaRVNBTfnrJdP+vgpzXHoDSYlGHLFG1tXcPxI
ZUy+zwioY3NbJmR/9AtJY+g2CiwdG1Qipfs8v9UTjX8nKQbwfLesohuOf3QJQ2E0
q/OQzEm+A0S2KIvUhSqS3fm/hutnWD6lGnk27nrzoCt9/zBXMjLb5x+0Bp7cE+Z/
UEVymPu3xmh+72XLHKP+o5WWxNpzFKcxM1iY+DdOWDH8IDrawmamOJvEAgnYW4Gm
1DW28AmzzZocjRTlBba58TDKR+pZL1sXXcIXzZI8PqXOLCtpJr0DZOXrJPrSzYxf
nqQUOR7jKR1kPbIiByCZUsiPi5QxQvt5E77eEqyLkoZEqIOUnhptZUM49kcEpJG3
DtNlzuSACaCxtjfwa2SDrO9GdhOENGIbz495Tg/fk9gMRr/vw0VE6zr18az2sEBK
SfGZRmye0iVNKsncFYSLV77stAnCq6qLYxBItglcmFg01UnhFbEQjp3iaFW9QQl8
LJgvcGYwZLa39hBnCKeb15MJ4kH2KwHRrgCv0SNa0UjrnTbNwKxSvyeylgvqRsYB
Zxl0hPY8ThScNA7upyh2lJai8eKx3TS3YZKnPpvWCE5yobb3N+/kbyMblx/ObNkt
A10n5t3dRJHk21eei7+K3OA0DulfZ3oerWps5wadkLc9PCmwaboZDnUqsEJZWyam
i+8RIIfgKUOo7D21uWjKW9YjXpq6sywhOXs+zYlBnA6lEz+wfcSlgHUfdzV1uPh6
IixsVLaCliFhpiTE2Zw9ciStr6MJQ7reCW5e6+jxVNXn3MOncc6fcZxNDP/I1Nzp
a/AOHq3P8BUk+IYLVyQHC7mGVT562CIcdJv+1d0cXJ7sV7VZs1bpUuP3tIn8NUMR
G669k0qgKqEdZe62aYOwvhAh/4oF02cy1C4AQAwAjYRCj6G6CLR1Jyd5+vu1ndlC
d7+sfiWWLPSQ87lqLorkPy3dEJlhUepWhAzmvUaoiEkG5hhj41W+/VUb7OYXdnbK
+Dv/Gj/NAUHyY2ZFbYBPdpdSoMjpAB8zowIcVg+Zu4noengn5ywSOjsdhwghUgbn
DkWTDiccn98e6S+WXwc0aM/H/ne+7LeccwQ61MogkQ/apU5dWezTNano/IjsLDmG
CFWWMg5wBVLr/EgplAvvZNVw6HGL7k7oFShsZEWzxQXPRwb2vp7YxgCuYNPxWrOK
I4x75ZMAFONr4kMZrK/UQY6XNooCA2XVKYXO91XXeZOXsKNidfaugv5D2zZ+i9rz
oum9M5WwK8wSgNMCreONdl1+VbON1DyS9QMZEmjFMNJKZls4E1ty9aI8nLNSfsQQ
8ugCGACC0li1nvo+j7/0BWWSATEbX7y/QPw1EOhCO1NtQgF3S/wpHFIYv3nrHB8N
cR7epjuQVaeVEdG0gZFnfUpqWsqeSZYFKlJfG8ylHHzNnwuOLye9B+daGLASyRcN
4eXpXNHoEpZK/52Bidxf/mHeOWcQTXvbqUVt5GtEUZjOMDAPfbI2p8YO/sfqgiEW
B3gLgAfB4S8RZGwsSHq7gAR3wE17LeJft+qHuKh/ZDiq1psoXuf9Ry+fOCn1EDUI
tk1zrDeGY4KDerr/8qu8PMyv6i8otS803KWXsQg01Jpu4BVy4KipJxNWo7Lj9Kvm
30gt5JjFU8TxtyVKNg2vhfsQC5pwBMvBQeI2+XPKtc+qu1Bbp3mpeBTyyNOP7Uei
1FHAG+8FZP9/AEMqFgFJJp0mQB6V/ZYOIUVghdgb0djHQhtRuQehrSgRa5SHrAIP
ZAp9pDwYhm5jRKleP/jrbwQlaUbGdiQqC75jJn5WM2uMzgPu1F0Xlp3yPySLB9OU
xPM2QWbQWTcekBsq+zTvIav5q6OroKdrnVeU6PrMTeK2z71d9Q5+zDP12+VqZIB3
Ml2kjleix6y86g5tshraDP8MBVoj6fJI+CwOF9EzyVtz4GR67vd40aHR/mwms1Xt
a4b72M3ECW9zbw6tit+byB62sBnRWJ/mVBOD+kUXPR5whlQvcBF3KWoFYFzEELwW
JRB+vE/PHmjP1P5rpygGo/9NueUK6RZQklJMj+tGAppeaBHNcy7lzLpGdArkzUoO
wmpmxt1yW2suiDGw/VafFKNNZBscWfsp8vFMAZJE3DrBGun2XV6y+TSst7m7NmKO
v16R+RI3hBPR6xjWOjjQckQBgXu065Ugg65q4mxNLmhQ/MYMTmN0V4rMEnpDNuX9
pVIKD8H0B0Au9tNjjAbHx/cbE1AISiFqap6Ge1DaLdQp0SFmmi6NitR93cIjYMja
dKP68mH61jpzuNz2Ec0Ng8RKaPzOIxwKWmd3DpRcH2YM4a0nPAeTPb/9J9LEXPYT
+hgfZjxEHAjRG8nN5CKysTegiD4yr7vYqJWaLfDxUqBrN1f9T9KQtMBvcEORRNNq
kT5Mug6V/fmNKv5ZgDpecjGRAQ+JJah4YMzw8irpAHRwX0dnYTTBpqVQVq2tUaHx
udB/c5nHGXUmwx+3Wcj6WWw6MCGocnozD/sTDmfFyzcxGe5B5ytjZBSJlvuXoVlQ
QEHB4bk+cm9whOmu7c7BuJPQUZB7G1cAS5SbsKeu1kiFheUPvXAZ09K31YgwAfqk
2pVKELFDYxVm8W6keB91fvv928c/TBluLdxuBW+GrSCY5TGFdYO2CYzANC6b7jj1
KaYNth7jJpr1CtpfeXFExEd6+4Hp6zFPGZrMs+MUQTHGqMe79q1ujuRRC962a6jK
+tJP6Q6YsuU/obRWXVnYOjQ9AxUCRrxcdEbGZ1cKRsrQ/GUYTON5ztBm069SdsAY
vfr53VdDEGrtHAVG8HZh1OFIm4gXu8bWbjMNVafV1+G/lVLz2+xG24rUynWiyxNJ
xOmoOfNbemI/OtmsgOiNjWLmW1DZdMXM/tA6zB9W8GSvThNLjDolkAaSp0RFULMj
GOnKYYdQF/zryvaORitRCRyn4Kgh35//fXHr9aQEkfc77S6btiUnzxFLexwlmqlc
Z3aVdmp779j/oUbicjk7Jsezo3ebDLCg+sIZQ99szdxGu0QfLCOfCWlMYACWIX0Z
fa7wMm3GJjMBl9crue6DNyxBxttlvjzGarR3wFzCMBTpzglvR8BizrnKxFimgBld
ypPztTNw+7kLqYM3ghVEdESkY3pd+uWM/ZJhiV+AI/fT8Mrkp6nCL1ADLbFmNV2h
pcj1NE60OGZDDiml3AzxW2DIdFGIIAC2dYXS+Kxycr1GjJ3huVWlm7O4pPPrMeH1
BpCiqwbZxRZtIBUKBu1EN/9HoSVPKM7wC0av7I1URycsdaCN+aJMA0S3TYZru0nL
BK+Mh3AISquHAWYWvL3CH76fc3oM6sXk8MQf9Lpj2jHlN7E3Ztyknbd74C+ljyFF
JoYEaTIePadKnCV+qTbULdD4AzvDjBVHa5XmJOn8Up6mqrZSNCqFGsjt2yPqlkmp
ncYvv245KV7pdzhy/PcZRuGO1Kfvd4UJbcj8lAo2Th1fSyaY+nxPB5l7s5K5Qmng
qQD5RbKBssJE+neTWjL/c2c6SJrQmIEQ6Z1KB8bsk6aa0L3eCkvvIFA1Ju0wsjK5
bvwBpdY6lpZbsWVKTLo2eKxa07h5wLYflfsmq93j87t05zLHLQ486h08UvXTTa5A
JI4Dj6kCwnRHlJqyB22WbKtCD/3uiaeUO7Ak0p7B1k3efaLd1vyOlsw8gNfiKLme
dK7KnohKI7yOkKrDlq38lxQZGdKUUVk8TeFo9vhFh5avP4K6uWCUGuUeDAeaJ7li
c6muwgfDl51ni4CLLvX6xu5FitabEi+/iP707XKMoiR3PhSDx1TWKtO+d7MOCBTv
VI75LugqkZKWSO85DRj2X+KOyqAVMWpFuUHzMgweRlVLlflBATvsDfh5cRP4onUZ
f39MnUtz4YnodT+sZaKoyLAPWjHIJaqj68yYHo+g6Y2ana0zt+dcMNNkvQsbenQ/
fzO14PblLDRzFDPCbN8R87m9+Tnu+45C5WU7Z1X1lU8QVMRclgOryIGg6/LNbfNF
ItQM6BStmEF7cV+x1iu34+GRoAckRKihfbYiGrcO2K3/g4upRM85tSFjHVfDTWaF
xllOKGcpEmR0cWpJDm1dVm0VvpQEHK8+IpQLbtDlG/lpGHkJ0qpEDZ656KaqIVXT
HtiTbWpesYWdeqcQiLopjEA3O2v8Q0ydSf7c5IFkiwBw2Rr350KCrodEhiQzTE8F
NOZHeiw/Xbkr0vMWBKbj34xBUxXTk1gOn3n0R4/OZK4R25szig6ryoRD51LrHl4H
HtpQ8G+9ZkQlC9TLRBWKXbZVlQWI0sqGxwZfDZK9+l77BhyWuLCjbvp/80iUop2p
a/hYjWA4zSIjeQ6GTa7m6c5u6H7n94z2f2ILk74aPrFHQOknTjx1bCEeCn/50RZ9
qwzcj2fWBX1glhQkBxzYQP1O3pVs6LFKIzEr6+K7c1WiSY6ZM+fNRmsW1pUnEJtS
A+CObJUMBi13eAyIMP7mJuv0pVtJuUC2dJtO8vy+feanAEoQQDnC81PgCeqgrhmr
tSOfIc9ENrFNZXwLI7i0y+32RZEjDZlk8P8EQVqUAmYoPHBSbzJwNGPZnvMKNcgo
s+vNrR5bD069JNa4UnvjcHkymqQHHHJZn2EGilQWTUVRdS/J3gvxXdvQ9Tc5FYDN
ELApnZ98/y+4RcsFSaMs69xxxGNGBv7gIQ0+YjdpKAVHsYl2sy+GJUTTBiy6lTS0
rHxqhpSfnkla6VTGRpBRuuyu6aFF64t/DFYnZOinwVcvta7K6PJ3fWslm2K0Cbek
OURVkaJ4NQh9WKwCl3hTEQVLQet0p7TYT5C5ep1C0r+VCjuhZRoKOkLAFok0hJWa
lCzGeoueJELyg4H2J1uqgxMHQoQBH5wV3qokv4ozP0VEWKhU6MpvihoD+9HKgf/j
N6JnvFIo8773DuPGHbx6XKoYEJXQGWcZRFkwc7FAq87tI/Q391TSbDYqQZW0TAlo
xKHtBLc7z8fhkk+5vPelo/zKXytlAth6ywpwIqIGBCrmp/PFOQRRVsRW5+ZRhfR1
p6JZ4LNU+JJDAjXnQqDgtfmTedkjEYt2wPXbQbbXl9SmOh7ojKq+GW7B5QGex4q/
1GJ1q/F4dyWS6Yo4UcOaDRHeQcSOiR2GVpM3djNWqAWDaePbdLByyTMD8FNYgLId
sb93EF9HrsYfUSCYHRNBPCzOmXpQ9KSPctTnS6pxVaWuPpyg+dkd35gWWkhYXgi1
yTRRwLmQp/A2rV4Hg98BHKzv3ksMpKGdaQ7AEjCI+KuiOLLFDPjfm80Yk+YORgjD
bT+5nuZlRoVcPBsHoJ3OC1SFY9Fpvq9gfcgzjK1Fm62/cnXIJet8mm9rkLBZ7v/N
+fgFWPV5Us7qp2oN5IjZ8gRsnq4dKlov3APcs6ZB6vsY9MB/F2srxri0ugadTkt/
bDT2DF0uIAmf8e4dn3Uha5L885nI5X0OaPqGY/Pjs0aYbHkOFAIr3RDs8FYWxioW
nBpNFMHmiKts31mJ3momgVZuDeMwXxHiHhgOg7gcSNqeBlFzpF6L2rUy55Wh8wsd
shcU99Z8KNlyAzu0a9qYfgw46E/QnxToOC+agVzAeVLuo8r/t39b2AsOc77xtlQY
bhV7AnWkCkNcuADZtIVdwpzxuM0oaoAg1doggemGT0gGzIy1E6e6j8v9AAtNX3F6
Uu7JkpqkhkOnbcMbV5dPZpHiCHtoA+U6X/ytiKHIGUxocZ7jmCkavRh36glY5Ovd
o7ylSRFhhz9/zTNBIlfbLyFmMrqXlGtCD8poA4Y2nyrsgZy6g//JCb7ReUuKjdyc
UCxcGtgDklHOcPfRkwzcCo/Vflf2FG7Cdm5X93XEXkjMOSeTV9S93loQ0D1RqRZ3
ckPoXBcksTUa0wPTKm/nDmIP6u99EaGKRbPMEM5EU8D3+tNbNDmvSlQALlnzYfTr
fpTGcotRIGTEGR2Xu80QtYATVSUoo1o4n2sF/UPhH747oduUFtMCAroR4tHk8P7V
NluCPcZPXDAP1zRtG7SVXgSob4lTVaVNfZyThIMPmCjYar3Wjayxz22ety3Dpt2N
vx7ut0RUoXyA8mOL7fTSouZaJT9UnRyM24mm4iGTtEHapyMdzx/XNBGqM2BHkW/s
FU1fA4oljkVvAsf0/lF3Ag0utiD9Ja34TiScAnOG+5BDgzWLaLsHQONairwdaPOA
OeBKIV5FZG/W1FwaXopnk6+KQhuF4v0ibQcby91v3JCO3QFiOSj4FmlZkhE1PTto
U4LEJ4cTq2aZw9Z7sHQ0Th61P+g70H7JuhOGpmYwyWTlFN0488CkFDR/joLt3FOq
8BAB5vK/HFpUXCb199ABZ/2FMq1qLDCqeyXv3dWz3dGyoBscGZeXqPMo9KVi/HIS
4oWohdanV2F8YVUVqxwAo+qBGc0Th8kGY2sFWtmCuEm8kG/g3KU7JCizWeKdlWFR
9c2iKPzbsBwnH9cN/VVsQecDZWnub8/UhMKdKrmUT42KIYinwEAAc6znFGTiyaJl
PuNcwIrt/QsJrw0cd6wnuTkjomLR/Nr9pV0JT0hAGceLOl+W7uSPHPoW6MjayJ6l
0q7Q+VSxtl2S7DPcBlGiu3TlfWQnu+EMz2Lpkm65bzjgufJDaR/s7z/iTDzP/h1F
2ExkAj1MzmwFPKy+3sOW80rfMe6gVrMf1yScmLbWcSTHvUHwzdOQC2nQCMCYE66/
DLTIL0uE7ULchjnA0eJbOfyCv3CKB5CSUzJuan2OsHVhh4jG2gd98+9aZvmCMpAY
2i9CeVq6ZP6aZcA4wnqKI4KnbUyu0AOss7ea0WcO30D1gIdSIIrA1iq/HJLMwTam
kWSewcYgO9ndNwnxOL+hrnS51cwxEFQEYxYk1ZmWD5AkZQ+iZZbkvOLExLrfiUwR
/gXQoW1APrlr4JzEUHKidYmYAucvR1l1P+SfhAcZFcRwSPQfooPMepspcRSbk2Fu
OreFvxvzq1Q4wiwDuon/6VHJTopim+ZNcgt1IWV1xHtwXx8IruNID/2U33IsGVT/
zzawP6td5yEaAvicPQJqkLIHld2N/s7FoL9m7cohi887ZNRX26GWXKNwKAMu5KZJ
S+DGRrZqLC+zwmX800PwatVjWX2ZAJ4DTsk4Ju/ONNaxY5uon02/cufATS36clBX
oHWqlN2E7R6hWkBE8DRKCdrPNu5TBnqU3rhC8W990YvOvDlOIy9p2bIUphwi5S0o
SpTyuNAYzTkECvHhKIOPwo4IhATgCM4+zDWhfvB57P1imkHMfYS0ltwBTjpC4eB/
FAUws1mwGK7f4ajtLtzor2GuICUXys6Y+DUJKFN8T/BD7if+dbSG0m7OqY1u9Zke
zwgW7ZYjO39UX8daiC4iKGM5eeOV0njxxwV9ocCJQJt1x0vFmSkdgYZ21t97yhEx
uai0FbC/NBPWeXGgubtXLj355VR4nF1glqXgs88/9nVoSr6SB70GmG9JF/3ATRhi
tNwINuNY95aaha2QZsAHEHRse7cuqfN7Xnk1GLd2Lb6Uka5GnZqOii2nLfYzW+PB
Xp4VFozAzVnPis9F6SpYmCQOY+ngEnXE+bM385i8p2i11fBsbh1ma/Ghkb3Aetm+
N+f8e4zZA9wA3/UGQrcAAvMy1fI8ryAFfdvU5O6MVHT3ck6p8u1d9/+APJ3G/8kG
2NgtsF3VpuTzC9m1xh7JoVJhwG3M6YDLNJ4hM7HYOIOYZxi+hnYnGqaij2s6fZnP
sb7zKdGwjZuofI8wbGbEvTasK/WXW/LYRe5iKpfFgmK/SOTxGUgIz7D+3NHmL3NV
VhRxwIPl8AI9I8Mr8XLQoCaxZe9L61g9+5JF4k4EjWIwr9iPjrebLu2X82kDy+n7
8t0xcMQzl+Jy8Naa5vtTuNlQUrGEu38VwwJzceyKxJH4NDsb59ZAMabbE/XIho3S
CWJG/QfDvWMqCnbfkOjkisbSEn0UG0wg+dRFyB5txfuwu4CEVt39MoCmTZxJ7LKT
4b9bXBZkRHLvQGx+gFVHjrFSvmyOGoV4RyGGwjaQnro5cneVKL8GtSsKIo+pacbK
OzZUdmP5AkhQtQpSlI2YlPBJwbiEawmIQQ3KCV394ExVvxj9EEpua1gy2SXgs06y
bM8AxrpxCPUMn6SL6zcMnmsxZUMArcsqj0da+tUfGmqDGg6ZDojQg1n7kDblmlAM
NaYRLjjz1qPTIHH/bdTbAy2ASOQdrls7hSbSmpVFsGd/dijUGUqk7Z1JCxFuTCla
Su2fivkfCYkkLQbJVAAJnZkmJT7YPJJn6yTecfKZb5KAxMhfK2p2NpB10awAQ0Lq
n4jzPjJq6F8Ymiv5TcwDM3dKFcawTBINyv5S4i7FsSsqs84PED8s4yPRaSeY5Pen
IcHZJbswcOgczXOKBX/ueYTdC2+Wbgw9GpialqUmXwkfidpVQC1KQ0u+iQUayj9s
oxVYA+c6i2JOfIFlaDh736F/1kGzuT+sm5hG708PDE0DUqaD4qukWjF4OYXsZFN9
BwCrRIxiIk9zWCWjctZtPOh2lcTp44U+es9iFtRBZhWH8GVUV5htFQgwHwqRQb6x
Ts97fAJ17lPtKI9ApAaV2fn5C/BZkgjnOq0r1VCdbHCJtMi+tEUNDk4/3J6Cle0M
bV+s4yBfbM97rfzi2KJtyPc05ndbEAZsvvFQbnJl22MqDuazrsEoawprGzrWx31Y
4TWopqk4jkZ/P82dHtClx+5V6B/+5eSVWujsuhkoP4g5Ou4DiW2EtK57iMIaGiP0
hOzPNmIW6wUTj7Lr+m6/UBvIC1kxVgavlwFSHBnsXVtbIVpraMOF/r72M1CecGw+
xqIKpbp0q7CSYyQ+eC5mDPi6W3zI8PLpkkQ/sMwy6bUkNkDbmjK5dpphsWEMocN6
jInb6YWY/98AOPprdRudgwC49jyEiw17J5u5qBHi51THjwhbsppKNE92TUdFJ21h
zQzZ9T+byjKEhQ8duaHQ7fMrP6FrW+kgbNlH+WWduZlkIO2+z1BfjhW6/CNLH9d2
h2SiSLjFK54tSbIpaYdTpxALZ1aaNRo4oUtxk7myAHPEVgLijHs+qFuTR6GJMciF
nrNmyh3qZI0UzXPEuINSXXvzWOr75iba6OFPyjd1MBjUf8vy9HGIspWpG3hxa4ZX
QXn0T9UJsRILGphXLHdcvLaSBYu3EDPQzPj9aXT2NVZpug+VrXQUwch/iMLpLWlv
Z5jKkKRGmqzM9243SYzYOMaEyR0TX9CgxSqqv7fPem21orH9e05iVFIFikb8rk+7
CdcczlWZ/8akwZ+XaLepgcyd53pZvV4XHe4qfmyZaKhvlMppsPD0cfDUZs/Wg6xt
GPxSqUmVi9ssQm0Zf2p3f7fj6ZQ+AoAw/AzUKUDge987YvanJoYFlZdn6A5FKUs1
i6aMmABYQKEzjF1u6yv/ezQcb7Q5claXRMVcwxXA99oLyZH95WEVyTn5tuRD1JD2
2QX7GRszawLgYXWGWhdPdNqIcKTlqaOQFei89zE7SwEYo7/wEonIAsvWyBBz0/SZ
WH0ySVB6EvboOdg7JyNMbLWF4eOjTwj1Am4Xr2zqW0XGTSRh2a9bC9NfMpgI/6YL
rPdRfhKDWn3Zz9cotFnXhcFq3bPnU2Mll5ZWaLEMcBda5m9skmJGETN489QKNrij
84syrUJw3K+qlysggbfsmq+RL9Mg6Mk3YdN1/LTO2f2Y2RjlAHbrB6Z6XKXPOkLA
qtbJGO0crpTKXtEjphpy5A5xI1br8UW+D2S7N2A7gJEgz13nbTRRPJiHkIH0fLxq
MAAjNIBS/+DLsFmG05wX+TyedG+1L1fiQOTnfSU6kbpfdYYG84H5JHW//tsaE84r
wK9krXvSa6sGolA372xeXc6x208xxnnh1UAbvb4C7Bnz196n3esDHTZgUY/cvDYr
Qed+kw6C0Rsdg+d/9x4W5qAS5vhb9d5VbgamD7HhV2VRj/Sn7sazl/o3xKKHbAbm
oS1Q7YJmu+xN8sEvpiFFuptUdlB1sBBXzstEKC+gSH1G8uGbgyRwrPKir35AIM9L
B82fHk0BNkv8VDQeY1rCGZRHCMdB448Yfe9P/V7XYrLS4aanR9vWq4M7r+QGYHFP
E7mhgOX+SgCQaPjMOn7n3HZoLlRwB3pSn35SC9y+p0Hc7x5Wuia5n0XESRETgXSQ
cxtGMFE9F3EQ4G7gmUH4am07oBT2GXhdbG/6vcaratfB/GNh3+DVgM2zIM5tlk4Z
e7VUGNnaq77e5uTAd7rPvQLlWiF0zisr8CcDEjreIz2kdLa016wbPPvrrRHMEmI/
7SE0ciHcnW92+PhhgNSmmfM7HIJ8m2YxkL4tGWbxkaZD/YwEmhfLTnaStdadL2J7
h2Q7ZlLCocUXfNT9dMQGEYd6eoC2SVBFokJDHkw4Nj6cMkPvcu//4gJn/5vRxWCB
c8a3GdJOU+RqbWesiAQLMhxld+yYpPyThi2Y2/aRNbZTGVps4gY8ym9tdu1vgUV4
PNXt63Srtwk1M+LSKevFZnkt9qhgBiKfyV703PMtkq97uKHddwbL0WcpXG3vGVU/
fwbTeN28lGvsCJvjygiVF4mtu6PV6eQDEiav+rMaaq0zSSAF0+64v+Miedow7bRR
JjbtlQxmd+btuBRmFhLPa5TA6YwD73wRNj0W2WOWHiVSkwAP4mOt5+HXI7s04law
Hi/QvmUGf3yMUDW14Y4IaE7zBwwYZAeQJyzAuiYX3a3ZXsNHDfLkC9TUaZ1585vn
dRxOguYc4SUo9/jPs3OtRjuaKd+0KEzrco02xssg8oIKFZcD8AANNtNauYnCUBG+
YKH2ECJZ6IgwlWstk8rTaAxJiHvYE6pGTO6JILMZsReaiK2O16F0DgqmkVh+f7oT
0yus6aJ2zNFFmf+JYuFQTiOCePqWgcWQjXmh2p+zOS0BNwFxi+TJIV6evdg5xA8D
lAVJsf8+LPmkULSuUpVjAYTAeQPKQKFJ8VI+UthuPCFBZJ9rpqI+GWf/BYB6XhjY
8hFeeRHfPlKYn3gSyFZ5uI1yVBtb9eRU39IfKI4Df8aUePnSIDQULumP2ql1zhvN
kktORfy27KM0cRKLyPMIH0+RkCbdwtEk2AaKgOcCtEibDhyc9iQuCllvQZ2SgPl0
S043Y18cZ8uGm/wiFW1JtTf4wn5IIMUDHIeQ/lWBOdZyqkqNcexGOamAVHq7vyMK
yNIjCmBC+8l2VL0Ix7YttOYrAMC8KZ5ZUTGxXaYegtA5cBJr/r4o0vYSD2LHSZLt
8JJXlt3DXsvuKG8qPkMRi4qlutGs1u1g/sGjzBPXcgSon+onsgER19wQ8l4sgi4P
P8HP/X4HoTZ9wGOcAhbyt8JVauw0gLZJzr9AULktY+0sBp0CSrSEc09hhzqrAY+z
Qta9SbuWSvIi4OBlJD48mtr2JOHMXsGl5i5YSO1kZEGQHB4SB4DLzANyLVWcRbE/
BIuqPPh82kq4alnzjwZ/ZcxRi+l99cqkEQiDOsAtNLPBruvBPqZ44oC/dJF4d4N4
cNBxUkIHX9ms4D1qNdr3H3dQJRWBA26pnydDkGb1XCWYtXU1iyI/tck2rK8MNdYc
p4ZCH+fgjMHwmZ106GrirIp/8OEwM6beQ9USAHbNA+qh3om7jeactUE/rEAtbo9f
9CLoI7RVm6dYAYLRrJW4eMco/a8OR+TN+2cjfeevOLlIv2gfJ5GBUx3RGlf+WyuA
M6arTnqFp9uGlXE/Qt6DJ+WmE80+QLIW3jPkaMzOP4evZjsp/1GNy7Xf+qnxCzbk
8yRlM0/Jx5YUgVRv9adjQnlcDxO9w7Wm42ZXU9gWTMdwrp8aUn+IJn1O2u9BeUjM
6WkNb3fb/h37MmuylrAQynGVv2Ht2UPpoYbAm5rEHV4IV40hbJG9bDwx8DQz70YR
poW4jtPxn3jPUzNX0RC2umhvMynHABC25yLyG5Q5F/RDDoUckJixTuMpMxTPRHQ0
irhwiPDbfemnqsFSp4cpbqLdFcPOpKbrJk1yQVac3fEo9tKMcFSTM15fICMBkrRC
MVzRMPTDn9ib1zxJILivDYhVvfpPCA2vNe6lnuPDNfNgrgRU0r1YwUn1cAM9KYhF
U+y1RxOLBt7lk0by+YhMGCqZI4yzG26imvKz1LlTj2lxUivnh0jslkjMsYe/Qog3
jHl0hAqtzjdKQq5+v0r2Z5TrlSdmpNSBVXT0pUcBTh6MbIJBid1eht4zJCLKw/oj
8lztYzcT1PQW4GRDJ90s+q0zV9rKW/cAABp9eOwVGaWr6CxrawSVvZT2swzuLOXp
pGFbyV301XE7MlHj7fZZU74dD/Eotxmh0s7KPeSH7M2kcQ7ZIVl32NXpIf9K4WPO
2cREgK5NfTG9ejY0EMZ+GTXhi3sIa6a+gPBVsXLqoWsdWR66sS4SRROERWIwmLFZ
6AHKWCzujinFM5SiP1V3RKgjyeb6xk1XYLFVNgP0HXW+KB9sg5oY8a368G0Arsfm
aD47heuqz2uJrzy1GtdkDpPG5QdLs0JS7ORjHaiSPS23jVpjzVaxpVww2LoohdkC
HhqbaFxC+TqUvN4ZAzs9nDMBMokez7XlaMIKHRUtmBN/uRr4XJ/mme+BXP6qHJJd
8GWe0PCu8sssz7Vt+4Kh8lG9pf8XKQBe/Gkfe96MSmQo3DrzlvyN/Wauk+eBlXgo
mF19gQMkhqUD3aCgXBhzpwzNNcruNDuRJcFES+wtaOae3qalqz+5dVyw+OPz/zJk
jej44uz6bbnkeTBAYwyaimIOuRX2bmRUjzCSq+AAt7pAibjU1efCh72t9fbdeZzz
ugxddOsUKZ1lW8Zn19oGAWecHkO4hsDQGMbZYfu9oW9OSzAO/yMQ7en4QfUoQZs7
/wHVD+Z4jzP418bDQiDw8Qr/zT7GgQ1lXeimuXNAtxF3n27+y5047tZVMx6BNuJx
2jyvWtSJTvDafowJu+wIOBJwUCDSCwQ72NyLm5NZww5+sim9CdpgmVoSsJ8KCoCx
YFT2o7H5dMZ4VwwC1vkr1FOEzIkOyYINNlFJ0oLTrw/8K61NVIWw0567TgTDgbY4
KuwXjIFTKA5s/fHr3wfOPJmrVv+LHrjGDjEy5pX+kdbKo56tdpRIW6vXam99LJFZ
zZ55B1qohpOHmn1tLWi3VbbaPGdJy/ilGUfCZz7YvJryzJME5lUdVKJ2ennagpbJ
IhXDQBvIdDMEvvaTb9foIlQyMz8d+srpx+trX1ptzf5ivyiV9UljnYfqiuraA1it
j9/i831iWn+aBHgDByuuJIeieZ5SgkW6+zD9gME1CCsHz7ib+46KbRaRV8wa3DTb
kItOTiPQKkOPf/1JPSVYHZz2vBExFqhbaYyclik2zljt6U4xLtVJ4AHIZy3wuKto
EzbLU1Q5N9P3HLVPZxWaf1s6L7YK4FMqXocjwHHlipDoA+a9uH2rD5zXNtSWFTz6
7JByhxynfjXTRX8tLiImpJ/wuU5g0gBa69OALI1XO8czVYoU1slsQ/0fjHiYs25S
vigqvKfwFVABV7aoHbPsHEiEpaSZO5GWnVQZDRV92EpQvQF4Hm6yF71VlRzZR9HS
bC26QpXwVG/mmTlAoEOpFAU9D2SZTdfA+wNOjvDXtkB0ostkO6eqkANBV9K35e1J
M/cxok9YjfdOlDQ/PDisS5G9gPpjuF9OD8UNIY+bWl2gVH5+CizU+emDjwg+HLqG
swQ7pk+mHgO838wpnksq3AYJY5kk98Qrj49EhoTXO2V/XTPIiCINgq++Y8hmz6Ox
jqzbejIutyg3Jh8LYAbxn+Sox+bm6qFlcuj+Liiipr3usu6/Bo/73uzk9L9fuRkX
86l4nPipyAIXutmkvryeQgIlj+WvHw5mOeB/01Xw3T2hyP4awIYxKLRipVQEK1rQ
TiLeZPxYgxuwPrqfRf/PvtF7PAzahN/iBC06ms7gJvG3x7SJIjVR18f9I7n7+wKz
vTPwfHozizu+UsSW+wcLv2y3u/uPo4xj2Jjpl7NP6qIt82pnW/BaykA4iPwGRJXv
OHZt6ruveSs/9zLUgVIPW/n7j3kFf/QGDxaF4WL8BQIb0AtIlR+7oEJfe6UIl9B8
+/6zBMXgRQcxuQI+9XRfOSYGBbsQtxSXmxFp4auxufLkFwU6DKy920sOLbqaJK+F
iH9p6nuW3tk1Gzd49dModJ+EEG+FDuetLPyI9eoi7bBk4qepKS7fNp5Pl7SlPS/h
u4biWSDulExo0cZ2nmChv2tVjpkpb6A1coo+P0QN9yxe4AjEVPWqDI5d3jiIICWE
gtSfFpm71pOmuQQRjV6gqg8yWHffQX7SYq+AkgJQJkUKTnMg+TsCGpHPUUWRsUyk
LZBQvUdS3io6vejmMOtIR5wydP8bMjyyttWwm0LAh+DPmOel3X8pB0M7k2z71V47
yVVQeNmHt0pmcggE32lz6iOscBM7CAACAhzgjykdb9pqzjDU9UpEtiDpgXmtdn5d
E/cr4qTBN3FJJv13v4aoJHFj8ZNB2q9q5TwwuVMVMJR67X47Wkc3XqEzMpqgztXR
umZghsb6OVzgt2kmzHsBMVpFOkNK2ocRsgW6sGdedmEdPLGe8DujYiQMflrPmRJu
Jspq2Nr0flp+l3N71qgSGalbrx6wGlWRfJJA7Q7OXwq6OMYsUqTzDqq9IPz3QhTD
vx/8ZnpTcIDhOEj9dnfWd7Q2duzrHCHpcAGJgp/Vq2uPsfZhu5fwh1LVqVCPSQHm
A4HjYtaVBC8rc7sMqbTNy8vdagkE5cefU2HHkk50JdQCvlHSpD+Nmkw6D84BdK12
BSZrdSXEAHa0CIbrQ2ih4Z/NZW1FDbglDfEbRT6xpD1x8OP3+PEPZZNoL2w0+OvC
7IQ72L5/bjuyIzKfU3GEmeYaN0pvx+Pe8RYPrzxUvIxtSHLV4+cO7eNhcONiP6MP
Ao5guCxwoCwKY4q5DRpJc3ETT6CiSd4HqZ/ps0ANLhpVER/DFEnNgSD14Ag4lW8L
8VMEMqKAHWgSG4TrgfkkPL9sH1criHL7EJiGsRV8VYoA6T8CfBaWps0zH9ahJxnu
7aCYbBaAinOkWFy7f+xrbSK8DhIhxEt+fTKYEqjeZ20kt14rU+OFrG3n/NyrTIF7
8TuWhRGVT6GJStgXxcpJ7h3dx8EF8oWCM8rHuG47vTfw+zQWX4L2JVSb3gmcs9fd
3OQMcAIHxCJ9/M9lDDXQNNaHjuJd4E0/TNQe9ulJK3Id6GYUCz0FUMXfQxKIpgYU
77tBHcbzZafSG+uJjInVqt4LsVUHA2G1b4jkf9YHzH3JTiYP6DGLor0uIJv0khVd
kNfpMeZSSSAW5mHNzVykVc3SDx4xmebB/nUXls+ZHPL/MWWV6ToTB5mGXz5cuLCM
TN/MMw9bzVO9me4S6JoG+jG//TRohpt4tLNLTQ1YOMwMN3FUM+Xp6s6fNB/JoCQt
gsFPXnkIWN55cNhg4viCs3/2I1S/2VlrVMwIYbnBScRn5kwWOEy2Bbe7HyfoFB3r
IfWtTBFDQJbwmEc03NhUs6YZGyCPZ7JjKNTi9oKNTkNgmsn8L8DFBVy9Rj066gBB
c5Bbts2/hHpUovKLe6exGVr9G26UMKPDPLqbG1uLITVhvAT83W4XFhzkvC/2KXsy
XtrkMWna2Y/mBN+SGl0gO6owufmKq7zhIz+LjPGwCia5EtZrl5x14NbJBfDtSdkn
y7ctVM/3xy9SBOXBjA38l51rmrUTGnzaSjgBb3Lo/RDSkW71syZ9HbJZt2HA5+JR
iSjN+0U/gQiwSSIAoNxpq9xqdaI/esac0+lJqWLjZJdLbnLMjqN4J72rNVyAUwM2
2EDtX32r+3YdzOuOTnG54r7TnFWRfiBGR+9LlH2nKfiE07y4rKGnYcyMvGEOLkVj
I80Yetqdjh1JdX8xrGqrc0HQG/SAWJb/UgDXxpTt3jnOc8lXRvMjkCCB1/5I2KKZ
o3sarXn+ZH419rCPAarRuoovNlLiYmKV5LXWObKIxsO65aDknAliR+/GhZv6Shnx
FDNvY/yx4ExAovdtJmzhWqc/jF9BWNaz4EyvjzlhpsooBUy5y8OBunEuskxclV1T
8mFEPgZcgZMqjsWbiziF8L0VOcDpoV/nhdT1vT3DqA60UQ7mGXFybnb7KVoc+bTe
TJA4OebIuMLMpJ6k/KNpkgqUHMjbJeYZbkq2XxKN2JSurU14O+wpi+ydkfWi82Gg
4/OpgZej9UiJBLKGnA2r2o4nloOVCpd0TN7JAWHjPtuwz8o4MUz5JmgiJ01vqrKB
+36pzRrspGtpQrBxi78PvkzHb6nJSKSbauLwHDwRorYEV+vtzwUpFgO3y+8WQ3CZ
MBw8kC7T2Z401fRzOuZoigpNMG5wd61cPaf4u3vZuQk2xbKE9KjvBnXyXM3YKMBP
G1xt83piw6Cb/CMtOOlb8gSOHx+ugs25hzD2xzUraFnkUEm7AYwDMKT7eD+hpR0F
BJrLZJJG/OtkaJGz018UmzqU23A29VzJ+aSUFxq/NdxcW37DhyeW8BpRWnLskgTF
2LpEN5RfsZciOiEgOyq9TnSnJYADGEvxgb8JeIhX50IoHzongKIAG5N2MYqYLlAw
90JemPTYDI8RE77R4qllomBcnXxbFTYLKPqGXBUiGbofADonnO9ECvGjrbZ9+uO/
xN7mHoXv2iwK6w2h3YX3V3x5xo8S+jHrX9rr33wsD5//WtJpZz9DtJV9g0sK/2+J
zn9s1A+fWupOA8M/M3pIqEIp468C6XJuX5p/4SA+4exZ/hVgY5PUxxbtI7jKANGz
kmA6aJ/fRn+2lgKdElFxDMqaCJF7IReOtoNvidlbPPkpXz0FapUGa2mSiNkTZTBX
voiRTG/cs6YZU4f+FCe9iZHPY8qnKwvBj6LtgJ6Ljqbjg43wMvT5WKtEuxeq7xgW
T6Dh44f58gZBlwRB0OcoMqS7HYTXcVwJHuylp9n4fNzcUDnLoYmRa6Hp1sNCIRi9
dNxOgJJidiKxvptXSTrjkhijGsUcYlPT94vKquGQOH45H0YQf+qWu0Z7LEwwk9Oc
ZsUhD0N9QK5I31PmXSLmZAyEe99YfstukUg9je/azMuPWtFRZ94foJBO7Y94YJIX
vw3bSXiEnHr2Mytl+dBv04GGWPTdWsIyX0gstW+/ztuYpKbag+gp8zljb4IAumlU
TYk81wtLipOeB1nhhUGtxZe/AhaTOm4PZ0zyMmfxNLOMoU6IFDViBt89LqtDaJw5
yMQaLO32Y4sOiGFsa6x9Lu1RpmG7ilo3giD1n1Dbd4zuTNyvby27RHXeTaeGRJsm
c4tRJZwYANWgTGDxgQvpj6Ghr6BL98IzqfbMHnoycKewttb9QoFkwNRE+aXXYvCE
WJGRUO96mQFphcHyL43OFS82OJ7Gm/cYe5bnTenHgrpaOyGjUaiihdobKhhfNTQh
D0l9TpzGSWa2Fgya5DfD+3xGnHQVscpCZawvST1+6mn3MN7uPPi+WxoFX1AgtAi7
I61RznmSMJrLxIFvbQKvSEGx9f4cjaHW19U8gEnsGhtZ2BGs0N1bBlNpGDN7DDgn
P5FW3QhC8hHGqvPVM9Hviqn2UQwVtLvv8Cf8Lmy9mS3osiJPme2WBv2EgvfiQiHJ
GkEL6wG9evljq+IYsjhNrJ9R1wHcVG81scbXnsyiO2D0AOHb6g+Q0gTB2GthQQIR
Q9/4P367uDZ35a9qIZlf+rQU/vUZWhIY6XsFE/qWzV2Ud6nJpBoE0a3hZ/xLWws8
1sv7CRVS2bQvJ9YevcKpVA14zqOLaHXz9tMI6waYlYregEAhwqGaeBTQY4TOhP/9
IWCcy2Kr9c90/zto8nGEgd5uTbAYnKQyIcJhsnYHIW5lUG9/JxjhLKtZMl43NO2F
yiN9Nx+Cp1IUvq2DKRZvDYEdrCGZp8ula2jtECPw0U4dqCiyIXrJMM5TljMcXF9M
BqpeOvF7TPDNJI2IfP0V5PvTM/sSayaa/b+IMA5g6l6vao1gi3ubjk/R5ZIdrnLr
LQ0T+Ib9nucU0puLTlSVFXOGsRxPHE0h5vuoSzv16Xopva5if/iXO8Bx4cQ3zKAk
fYe0ELdJErioXPAJGpk81EaSTLbwmSVanJ45wOUwuFLq5Xs9r9SLQHMyT//u14gc
we4H3mfAKivThjq1Nx3h1FO2V1BKyk68xiPqnMOd6mDEKgL5N9LzZDuGsJwnJ3Og
5YaJQ7sNacLuSc5WKENzhpACvs0Hr/OC6qSS0ktJ4G+8zLIMUUVgqxpoiI5XmbDg
7AfQgRVlL3oGyksgvK3T4wpiHa84RGjVxlVFXrPcWezvsuKN4lP3Mf+fwHvsSw0a
NNVMiuTt6gdGbulL8/2GdyrJZ5Yy8xCHuhjU7ay8pftruHDMiLwN+SdRSd4/DXfV
vHWyNvOevTzZM9xoCBx7YKgi5NxRp2rfcbeKV/gCGSiy3AXV7d1YjCjfqnnHlW9r
OjxkPfcLuipisUcgrydDCP7Y2W8791XtUSbs2IZ7K+y9rXmC/CMMYAUHHvCZCdoK
eVZc6+zXACHhtvOyQuUJvz+RntKdFLy4M3k6XYeWqEf9bghkvoawO5P1vIasKLfX
Q2TRbudE2P3k5j/cCIe0nPj5mapqtscD2UOGHCXw/NRgyVCd0vIYgEZDIArVdGT8
emzKOIBli0lHWxJ+dqFtMmzzGBArm2BFXJ5QAH15x1dtQk6R/q2NEIRlVeYLyexN
HsU3d1q3maj+U+P5hu8AGVCFd0+TKd1kiTXx4Trh1vdJPuoFIQSuYxgd+1sSU4Ia
Nj6TZ5XRQpGFj56HPtA4U1gTrhpi+iCBi5SQZlebIdUNxcsAtZXNVW6Qr7M7FPB4
dxwk8gqNB5lQeTNSXrfkQoir61Z0Cgd8tHuAzIuP9tsvDVAD+LIFKt/aaJ+/XEnk
bkUhNWU5U9A4/XOvcEtiuo8javQmANNhIH71W6VXm2jkTN2W8mxYJPZiC6aC3Pxv
9S5Hl+kzydkjPGJKeuvKzU/nlwx8V+5H5dQ5jvIoLQsu8bDhiB2nwBVw/AKHrz8K
kOsx7MBqYt4v9ipq1lL8YFEi5YcuQXW84XaHsS+xUoEe60LDZGT5tAdD6w4tepEy
7LCbddStbIL1muzrQem0WMT2rtUjJa686CEe/XhXCAIY9GLrMa/dg1lY21+a553R
VctSGQ4BZwZHcrNc9tQnK2RlCWojIXRC1i70U1L/ozlkN7R0u2YrPobgXoyFQTE2
od4SBpnPMWvMTWBp9Xko5pWmqhCnNdk7S68Rvx9S2srL2aTSFj+tHKE3tPUFyIN4
MFq8GGWeYv/hSEIyqBl3DHyzC4Xt13LI7cZMYoY2q5kBGr9NaRIS4YHIqy5noxg4
6EzlEIiVpbczbx/umEmHCRK+D6+50/shHt6NUIzJ4Ts4y6bqik9P4t3i9zvrU1Yi
qHtph3d+Dnj1I8dqEo/ZhN9HaHt1XI4MqCdQ15+P6wrHsLa5uruU7HLUSgDVeuxA
6CdxEVfbqMUawYy1k69CoB0fO69azEGdXQ6TkN7vDReZo1mmiI3MBA9IHpZNaDFt
yJ9c3yD0+0mMdCfkUCZ0ih6YZgCvWXcXvuJGxThLc76lJ0v1/QYckzniqYLVxiXW
aGwhBThBqKiM4J8bY0CKuKzlpAI839mm84Fv8AADY8BaCvlmK9H7fJLU3OXO/ugY
7jUTKSjqE1SqOP8W1JIauSjr9BLbVmJSu9NvmvtDZANakOR0nmmbxWi8mySm6aHh
6e9lrI+13WgXgI6+5MswnjqE1fYARq2QSL3wl8XoQxn82i85bRWVHwM1bW/ZaOdZ
rI4lrfMhk1TpadgH6biNK9MLVziVZfawVrsb8tNu6LH0weqVLgUIE7519vFZg+xv
vSPIEBN0lIjvCQj6a9zUT1ZHGkN+0YMUhnwDpPRhdhJ1jmtBs2Oe2Grk92/Gn/jU
PYeAKwqnUZdD5kYZYcQWusSPVL84J2YOv4nU9L/Gv/62vWgi2g1ts4XX6/mOMXI9
//4svLp0GHdWv2b8/OLa/fyvwOJ7aYCvFN0vT9PGShc59OZTZ1+oqRKfC+IeX99K
Zw1Ffwi0ljaUpcmUe3qxXnutlb5+13l5qOBA0ZuyPUpbx38RsheNPYLrIeN7cOUg
qAmx83NKaJ26tMVcz7wY/X+7jQ8LjdYxfFu/UwhwS2ggTNrrtI81FVzVRlBjooJf
2yNx/P8mQWrJ9Q5yWBwSytGc9nNq+v7NTNMA1O2dq09peZIjrdB3QL01BEMs4HrD
IKN+oJAeNKAWmc01J2zrAfKCYDoJHZZYGiBrwmGMWJKxsGIWbuWLGpInh5zmTa/Y
GR2SAtUZjQDzO0nTmxIbTwgXgi+xh0YZtC0m/g7p+zmfxWFfgKufQrfXe1duF6Ze
ofy8d5L122UZY4+oKhpVyOzBf4JmRdoGQQYMuVeCrxIEKV7QFNPPkkkHB++82XRk
yZyEQCPH8pDnuJHKBfy4x9WPzLtiYXkZQ1oqhULMDm0OmQ/YddtX2FngnvdBAK++
sbgh9sbU/1AejIUIe0YJdLQKUJd2TKrH5v0PvFB9Ko+N7WAGnWwGBQjrq2sw4VMf
M9b7C+nHqRp4P14MlmGMO9m79FNQa4JY3EWQmyYpO9CFpwVSrCSbqkU/bA/60EZ9
YQunrwLnbYXfkKl6NIG8tkI4+jIo0VhW7tHvHT0X4f0Qr+8+aM1Rn4Zcv20XqGZp
JzIh4Rb/gBa/atjb35z/nEaEPC7P1mrOw8LG4xb63P9l/bwoO5PkoxKFidX243D/
CsnXOXpkergHB0x2juqW6mavgVl90RrCGIbOBbsWHhfWVMbfWubD/nNtUS1cfFGy
oFelpwV9gzgmnuxinvYw2AHlA1xsgKoVMuG5EeHOOf2QPoc0Kf30QuoW5yp8LB1g
SKIk4CDZglgSsMrU0GygIGdqsq5srsuvQc7vPM+i0YqL3zmjRFSvkYxCJqIbeC7p
GfvsBq1AEpJJXqcTHIEgxaD+rkqlohfLGnfKCoK9lxxBIT4IVrRYUPk5/7pZ9sYu
LeX/cO72Bmv0uQPclu7r0ZiRaLTpwIrBa/ScaY3JLRJz1fYnsKKEieW6McM4WkZn
ex+g8pdGeZk6Q5iPZfeUGJ++t/TCfoPpb9QH/BZ+WbZ8Yw4MOh+0B/eZZtS/kw35
esx3cDPK+cnN3SPM8c+Vb0QVbXcLUbOUTLOpYl/TJY06rjCVYoC/dlsKnqAceXfC
5oFn4AFRjBwAe2HCdaEcEBOIirxkTmyo20KkwMmGxZahU7j6e3wr04UKmWr5eg9v
kwLmBoz2XHiqej4C8aTMb2DS8FZocfqcxm6Bst3d3FQfpKveWyE86AAZ41oqNhhG
yJaz81XiKeQ7NefJsE4omzCPRIey0ijXS/hO4ks1p1m6PlGgRUqxXIeJZNd06jEY
z3JqUkqLKj2bLCjvLpxSxsXmpyS/hfzj3dwNGqqRDDhZl7DfI/9wFTIVLx9zBrA8
DvAo0PJNDzuxm1q9VhH28LbZIgdC/KWDsSeLYTNcBaNJjx9YRjgNu1tcPDalvAXx
a86YK7LRjXe2Bgi1S1hvEU7wI+GHrFdNOtaSmvrhojRAWCI9Jb7uoPj5NQN+H9Aw
nKqfJ2iw0qolNyfFg9DnXva3h8TOgkehW8wEAEMch2JEr6Iwcj5GKREyLTeA6Ef4
2ReRr/c27BD87pBtZTJYkTO0rgN1iujarirDiozxr0H+5GMStbN0ZwP/PRCMMLuJ
z2WenkD5/UPU5Evjfj9phxs4LmroE8oQFlwlPYDBWkt09eJyl4yItFBxR+5yTrcV
VIMa48GamdytPIIewr9NLEKyfxKCpJ8pLItEEIt+skQjZLFhG3G+2XRhXYdsm6MF
vetpnHRTh2O9agWJdJ3X7F+k+OQX17lyeqydt0HHvuwOWBWNeQ8qzN2+ya6Hte/A
k4NqhisOxc9tTTyf5Jc4QkO+TfnGz3Z4WQLpr3qMHfm3XLpGgZgnlwDRgaz3+Wxb
7owsJOQXrk4eKPEw9tM/XOci2VFO/CPiFcpKrW9kuksNGYRojEp3sKMUMnLYSBjF
hY/vNYevJmLiitk9kUL/kAHAqgd/+eRM6pHibHBXVVJBLYgk0FwFlAXUWZmKUuG/
yIBtnTQSPSXXfgWAV5NlkBYNEj5br0eub/yZ/LmsgrRC9zJqtci66UcteAOAmM5k
ojloAPhRbEp8aU4ll1lBVzcd86beY9FIo9R+WSTN/rjFNfYu7c0IZGj+RjkkTn53
8xDsFiiUm3J6gbxCDkjH7R6iKFowfmr9kbezHufOSv11k5YaW5UcYnb5ba0dqYgL
+dUR4yxdrcQCQH+/8vUrfrV68wdU/K8fAOf0n6eqMqdwBOc/VFxIfnca3dDPMLpb
pjyuwsJK1n2HbvqOfzoXwO5yAX/QQGdejyDdsnf3/8cIkQcRBYxUawywoE5fHr2Y
u+8xO9lCyN+1zEjHI6Kyw5wyp07xUxTYt+7P7VdIU0dVIp5c463PM318PKDFRHRb
3+E8naZkJDFDLDfqM/mMQ1unGGHPoGeczaMpmMg9IUUHtV/AMB3oBLKpDC8oM4Jj
MoiQt/6se1PUgz+9KDKI9qfj4xgNhemkeavMNUHF0mZpTNdIhV26npKkmUg0XuVk
zAHI4rY+L3x00LXIDBXmGRPYOtmP8JOkJMfEn8XUUMxaknaruTOelUKlVvuC0XI/
QheSPeYnEgXnEqHCpCgjxXsQ1P95NO13rkwPKvNHWf7iMopv5Uuc9CX28yS1u/FQ
dkjRniCW+l+FqCRzEANeg7sgcpqGRIxPAeE5JO7fp8zl+7WzhL7ozQhkSHiy4Ci9
ZICTDMo+1RTfznpXLd+9EQIkdfxshJemjbYYfpNzLZUOBKPlL2NBeNOdlIG9az0i
dKsquDukWCS92u3B38oWmzVEcW7RZ+YpKWN5M3pkdXjwkchcm/k3HBvI7/NZT7xD
/q6ycF1PwFH9tN3x9h96yzlgwLgx2ypaKjJ+0ZXhSATfRW2wnDvpm2Oxkt23d2zA
rKEt2+z1tCiR1KtBnaoHAv5jAgK6qfGAO05fpYLWjEZCgH2wLG1RJpK+/t+ZQGrZ
zSalu/2D0MV6wyQHJjoQsIHJBV9AwUp3oxKmNOURGcNdprSK025Aaf4KmsPlH7Jc
wdIKv4BjkzcgUlTaAFr5mLTuT6aHuZ+BQiIhFV750dEYKYPtMaoQ/63FDzogokfF
k/EVxpX8sP6HlDdc9WXAwNRiCd2ZzF8hP0hcUC+vk9d4IrlHSkTSWKyWnLHe6uys
q0KwyRuyaGHm5sCBF7PGzL1/QT/OO08fU/a08v9yj+8ll37ZCqHBiUzH/bdOGHdB
O+LUgzhCi2/KSFTsId/vO08GohuP7zQLh2xd6GV2IcxzUMCmiReqF/gnEuNk7BHS
OsmlUCDx+sfA3mH39jdfUxF1OEcP1hxpSZDujtgW6ial1FzYHvQnRUeDeP+mEzYQ
q4YWl62eKLZT+kCzVrD9iz2hYAc75snb2Cxz1+/OxzYuXZ6vX+KDlOfo7u/mah2y
r5Rt7pKThs95wc4wnelqfwP2GBdCz83O5b2Gr/alkuWiXFKsPHIOz15TM5b2Ff5v
zIQ/EgHg0S7+CLGTV8Vo0y67DAt3T/NUcvap4SorYCIMMOmS5pFtY8IuwLMjaAjj
kuT6rMGEjTRXLy/VghJbdn3TZUm4+BlYHHPpHtubXlLM5x0e1WKEhRqNsr+qXbOh
4Tc5XNvyTQu1LHAYcQ5p+Ip1OYSIxA5ETeTFLs2kCvdIGw6NY5vDysTR0f1axYUd
Koqj/hKgZTZ5W9clk268hMhnp54a4t7qRmw0V6M49xOv50wjVF0ibOh291ZUt8nG
x1ll25oFfjdrtOPCeBjbZ32Zg3CNIb88WOMqNyJ6EHm2OYdkhCLeCVpdRxVcHcFS
x4UKqWVOfDHht8z7McWRm7J4w9Sl5awrHYVfy5hAZ+zkr9G2UyqxhhY532zanmoK
3ZbC82fcnu5objh3SaPlBsuHBLlnP/vtdOfvyU+nlizOwO0ibc9+Tc2NWk1ZsWaX
Do6Ys1INyx6F7H/Tb3QPgMcoQkvYIauziqx8ZHdmA3WQsoAIDLgDewZ0seOCNCAx
6+TakeRokGhBdqIBQCjHBklsnAjowzyXgkCOcJTRsuDkJnOymYbQahdgboi9Z8xD
ItgDAnf/QA4aFD/59mninDSgTFZ7coqCpUD7hb1ZDAJM+RfxGU61ovtf/t8bCVy7
jdCbeAcWCWU1zp4YfimTEUJpZR4NI9KBRNkpvKJvPcXcDy4hO8py1BqDOBy3JBsD
+CA9uPVedvJ7qZosktlZrweQyCXQ4/TtIacp0ShiwQRpuw3aqC9zaA7BsBKxfhp1
7pFzFq1FI7Lw9WJvLtIbX09CZn6/RByIwKkSk4QgKClXfl86bZuHOh77wK7QYJgL
q3WzIaWRTPTQ5f0hvIVotniJ3UQU65VDU8P0l4qZEC+VHo1ikHJHEfiGrETq+y0E
Y1Yap6i7qEq5hbtk2HpuxLpqMWlr7jAj1mfvaMRgaoo+w26Qxvw3yJChuurIh686
94bnj7kE4sO+yKiGALvSrB6KMvlA5gsYrn4adJUlKrdlHjwFHpE0aawmY8OuB3/P
F9HNxpHvQrLEF5GQufu7PRM9Hit1PV8H420HNeK2Mwdf13lEv0QJ6QMv3faiJm6o
SnutxdBxUFUkCYSEbqCIfBxY2iGvAyebM0N7BtttVmBaNqIH9RPdkhUzDdVCsXuz
9Y0OIMGmvoemRatgnDm6LCXr6bk+ZmaTs332Qe9MtJjk3Hq49+w0iWP6ew1MSr3V
ABl9QVU/Hf2FP4qWk4VVEsldabQpDKb9+rHH3bY8g6lEpHaUqeDXuhUb2vuMig/U
tuUtSu0blCG49ENT1mQAKq0WcvDPw90VcLUrFS8ik2MKsufiRYs2zEIpi8+vInCk
WzJu/WQFDdtvb1PwDSzNUymsgeMksdK+VecRv2AO/hGu2YhrmVz1sAJ18U8EmjdQ
B4P9wmhYVzUIuUdUvsfUS7Xo5HJ2ADyTmeQjx9ECdhXrEInVuZeK6kmVwbm9iU7K
/c9w4DIGTJVSNT1sLdmwNvJZzwF75zDr8Gda1YrYqbdXgZ4jpuoaupaW8NUvesgt
5gWxXcE1k+v6sM/9hUL8HICZkQqzYVnlGVdVfqpe/g6rkM0g6kPE5qLJAHwO/lgR
oqGF81d7DadlfDnzY2gyVKkKleVzkInJ4u5+G0DL6fQMkZEBah9j/7kqILveOhmy
38tW1EMUVc3BcootLQzZk0ZU59b2hl+LuDV8YWjveNWtKMrpy+0PXbQpkxXM2fqH
UXTJU0gyXGgd0TGvYH4pSVIJGuWJbtmvj2Qnagl7HIttOfBe7AdyCc0MmBFGalEj
rkqi424SLwCPEWg+/UsGfbHlD7FFYl6KJrhHDUnGXo6eIG1+OuGKJG8CrdVPY3Yv
7mMPPagrdSfruNhRugUOhgJgXRB7v314LxeP/tW5/amYVz5LLff0tyEkyxSzVW9Q
CPxhZil30GOdZ16NAP1do6FG2mm//7Ka67g9zmm+o4rNcpA5KS7rfZxP3jg5IaEI
p8Hm8gKhTKaKh4ULD4l/yb38u74r2k17Ef/i09TVKOEEYm/MqtpN4V9qCb0ecVDQ
Oqpi95zRTLwNhReH7UQUsc3BC/tIAgTL/6UtftSykcoyCT+T3GDnBWew/Hh9/Fkl
3hRMVImyjTh0eioqjVt51HX/pV51VduZejSbJ8mDgxNwnJUlRQKFlhKP8qMUpEWp
MP5zeEZ4QjTsLnwewNFHW7xpfc/xxs4QlZSM0wwTjszFnAcGDahtVmtmIntzhMXz
nOTbSVWJMXr4kSLJORjv/cfXKbs5zoPLzg08aJ8i8eJ9KNUnsdjc4f0QZlZc72Yq
6pK0i2B1MR27PRep0lhRMS5IjGFbJ/huoz0xuqT1XuVABA/y7aKN1/QN6mLaqWNl
ZnftwiDnxMYmUxx6nw7pCFsi3FOFkF3koSSHAEcmGIdYwsehC/1zsGxTd2fi7AoW
vx+5puPo1to4Gsx2ncW8Z2n0/eR/vurRNRkh5A2MLlSQKrYUtgB99bCITNCb3Lju
CDnZOeargkmYldqlM091pkTB2o0CZi5TSQoifU1gEU89LvbbRKcLQOyDIONfvOHR
2H8M1umMJP9wYgqkw5wtUOiqUeQqs/rpkcal54lFbUHX6KYTHsf18dqtpLUZHmcT
hsO2r+cW9HHF6mmH0DYntVM7P8MRmf0w0BZywp6zhKUWUG+c288CH8sIpwr1whkS
RB6w9FHBCOs/Ew5lnd2JN/cph8plTC8GjBK37UgS+7+RT1S1yGb37Pp2E72KvWmI
6+heFyQINtvYNH0jI/U3hJhR7nZFyJZil5yc6lHH+imnWLClJjIrjcnwQisyQrTH
T1fe1ygKKYYqRk97MFx45o3Nf/sEnZPeLmRRTa9eeMxXNmIAShj2ozjPZg2gEVAL
3VhuBqKZ91GcNtIU25FDppn/McLSP+7/Bm9S8RsIQg/7R1ANuzOKq2YNgmGev3dd
GYN6r86/3h3PxNWHGa+apXmO9QzWmBqhhCm2bC/GzXoNWqSqxOc3lRzqrCmWbqyE
VHpZ9tBH583AKWeUGRZGrTH9eMLBs059Y1avqb2+HkhV07dPY/7R3UKj7S5gtNcA
anT2AbiJbzChs3sbftUtvAEJ1ot8+mFgT93xstM2rxkpKgpnUJ6JJFflcxbNd5LX
RHl3sQJ8KvTTULXa/WArqI1CIw1eyzFYh7XIBoapIOTQ2/GaWsculsaBQD1jsMRH
T5mSLLZaGx3FHO60DvYfoajDq3OF4NsHm8kzAqjZ+9ek1eTY7FrNsG87BW2tWPy5
tkvsV4d5oOQltnPt46Xqw+u+9d+Ujg4VQX4QsoCNl6K/5R+/lM0bercx0DRiBnjK
wau9B9FjZ9IpxYS2/cKWJ7tYxdJ5pduCKwF3tFC0erGiUDHLkJU2MIIqtl8gc4A1
gLCnNlr0r9bOnqSb6dbQ+qMihmS/5I4j4ED1qS3oA+G5JuMyTRkArDRqJY+cJvwR
cokK03oJqAEMnnwmcQwOAyucEgAn/7DRSRRUPVENXjztblTQliBP8dIk+5YKPl1g
80wFEiulqZVgSme+KgKeu+v7PmIiO1FhH9kIUXkxnoAYW8fPg9HMW698R0rVee4r
ctmog4zilyqPM0xykOG8msLSH6y+eBy6rHDCyraYkXz6vUExP70pTjeHqXqWrNni
BD5rNPEEuPCOFiFMEyOZtBd4hppw8pwHzmjgAV//+46Yrm2cje/+8ACh2MsWg7R/
FxS7Xmk9VrcjrNNzPvgZFtdSXZmU6gocnhcQlw7CeXafJzesouFo9ZZJXfF7K2M2
1EQ9Z2wGiz0bnC+9rV/LMyznVCfk3vEn0gF/F899bueDDXO47csTfEEJIwnYBLlO
TOmOqYwqaislMdSCs+779ODlO/YpQqk4A9StnKTBSGp2dHVy7r1C7qKgCZBrxPdK
MxJydH2k6EHu5tdj8m0lZZJVxXO28+DPc3914WbL3lJq6CohmcMlWy20lphGj3rY
6bLX+kH6yVck6p8HjnxBROFh1JyA4JkwTyrzBOGGKHCIKsA5/X5FV09YR8/puQAA
FlPbCysc+mXLkv+7JNrgZaMwtebKG4HtqK67PwRgFalk+nEuX/zlp9KQ2EKzW7SG
gtQgzD4pi3nwEB7bRg0HJkDXNkx/d/5mUJK0ZECXxf2mIjcqMoxZDdCx6dLvFz8H
RtEngNvZBBF2AYD1phbXZPD96xClLeG+wpoC3fYC15ZoYHUca+E9M4GpWymR4tFQ
G0OY0Zi6HdVA9WFSua78TbRwXPjaQBuZBmrqVRf0H9W/aUQHNvSWp09Ou18xyMmh
I16RyA8YijW7Wf7tLKIbgunqOKjofu0OK0rLl3p30foncL9GdJB7u0lZM0RY5sk+
F+lhQ4stC2tghGFG2bDOf6mKBTmGL0D+dwVBzebHS+Zmf+F84ZMX8L5BidkooHaq
INVZzkBUhKmEowezGx+vM5UAtAjuFUVDfAsXqB5T62Rl8goMaGjnTRmQruaZ24Vb
S3dzYxLU2NPgqqA3F1u3TgpMwW0z8ZJFO7LQ4hdhTP3z4QAxHGce8Gv7NrP7eXZ6
kTwghubrCNjtO7g/t1QBRZOiHmdu1X2ePq9ZJ4dG4kvjhU2jzf+AE74gk41jztvR
gzZbJUPNaKs+Iv73qXRiXjDL4ktxG04reXy7ZgFHqfLarsWt0gMzhS+IIUwxMSsh
bE/6XLN1/MsiL4T04FqZjEZ3qwV+hyuzqwM/H+zkrhLccfAj+078alf/B/Bem+Pj
mMMtIofGXDAKfbGpLa1hjpJYxue1U6h/gOrOPOkd37pvZd7cJ5R+1LHktEnT75I1
v8V19QPB+EX8Ar5pbM/8asAcXO694j+Gun+KVOCtWLVhb8qefrKp4zsMECgPE0ip
2v1dBl9xXKlDvNG3og5sOtQDhm2yl+VEC92giw5qcvvLHO4By3GlUbLmGHeubovL
POs8H9Fq8zMiWcbCCYySA/mUytPtGxexLw/BH9ySn8RMrLSuSlfbOYDqpb2N2Q5S
iujw6WEHORGfABe7NireakVLm4LV73XOPv0SOl+x6+lSTR5udCZF7KuRTwzKpOfa
Q9ydYPYYaLnLWfhQ3pNR1X37FEGl7Qch8klbEzigCGDVPEt0HQNepYXO0wMOYy8q
6ExAeotNHxktZKnxfM3N2OXvoEZHQcVKrA0Y6CzVMGPngwwd0KkjMUyyGBHmjK0c
kP31psfGjp2rA5SN3xGrCE6hLoZ4HTtXC/6GuduKtVaRfzt0CD24qjxAXpQnxTwm
RmoZICwdMNvMFd9g14BxU6r3IY7KGxKePL9+7voHC+eaAI7m8TgYWJDiNM+yuRms
Q3yMJAs58ZU50eT0bVEe/VPwF4Xi720FFxPZ6X4/ehEVwsI3D9qTcQbruz9uVH5I
LxhIg2I1B42YOOhxvUk2lIKVKwPxSD5ATKgZjSkKUtKBW4ra18+X45s/JsiAOP49
6vbzGyf7+cR5Vm701IcgqW/5o/9Z8qwSJrTyvARBanpbds5gSw+ot0ZdqhFRnzvb
d1l1JAQgbySkLvpA2CqWF4IgOdvmiuldSxQvoNMWRG5lq0yJ3Rr3hxD2EWTtpnR0
FxPd5IhNKvNJV4skmrdXoD+XdM5LSWmrYtH35Cos0cuCde8E/KBc1yienlsVoOYf
6vtE+ylic/hopwuQut9QHysZmh6xrZHiQoxBuElv7A6F/ntWdMLCjVCmQl4j/vO1
w8xxmMY9oIM10Ml0MlQEEm0r+G8+eGJDkzwMHka+RkHWNWB9JocD8uJsCqORPdUj
3zmH5bQcAbRRkU8hLoJJCfQbec6IRgQfZ8lSwNeUL0lg5/N/M6ynqljxENpuzwTZ
J+HcJwHPpmB86FXJIqKgnnFVEi3IbOxUMAXGQqeG098H2pphNTosIWqpyzZo//wA
iLgtfpNlEUueuLuQrvOgwL+XY12oZGUIJkNpnG+AGXUxRfoLaxZL6inNGMOzGUMf
3068jkXdJpsd0dbr/xRWhYebcaDiZtetbc8JpxeMtN+OIiF3KXCbsAWGXgqHNkUb
ZbqO4FXOHEZWMtAumzMK+s1FJ9VJ868kAPPG3E3Pk2XsQoVrqSwp4z+Gji8nsg5M
eY9bujoXVzuCFwS/I9TExWJlcTPpkPt+xWIeTPn1lqw0RYOZjYqp3Jn1BLoxjexA
iTA/C2QpHxEcXdCI82GYACtbdbm2dHFMoJ5vqN4B7D5eYFZ115bxDjZjwcXHny1l
GEKPWfZkyz0BFYy3YDyoE10DvdULtxtJ2f2sYM7GGeRTTxfb6SIaj5Rm0Hdi/xxk
KQCkhN8+MlbNWuOcmJOkSWqE+tLdoneMGUFPqxPe9Pg8PgYhj0U+qwhDC7s9P5q9
44ZDZWcGwFqZhcvtzhLXuQRyWOVIye9SDZe5523+hYiezLV9bJp+mqkdfXWmbUbN
LPn7wrp/3QvSVoSzAol57Q556xKoHl6ziEWhGlB6ZiO6rr2OFX7Zb510syNhVNwZ
rlg2ieNvmgoANXQbsJJ9WUk7YXrKwCx9nnvtiG5g9cuy8KwdnrQmInL9Wub9cUKF
4y+96Nc964Qf6q5g6liJ1KtBy7v5ym/Wn4CrMSoIYDqeU3ekmGvT6qEywPlNDX02
nhT4Dr9YGDsaK7eMZuRmfy8GavjiqRXvl387qVre4Lda3MEjOGp3+Eht/1r0Zhge
ejckQGOYdRHX8DePVpLHf3Y5UDdBHxbVIFNGbphiNr7GQjLT9EUGaUvaSdcEFgUQ
FcykDcp+b1BR594kHBTvgMiA7q4fNR5OeFZYE3FRuKlEGWnD3dkHOvrwlV4vqsq8
3Iei9v8xhM6Mef07utUhLI9gi5/e81Iloole73HMfP4Kz68ea1T/OCo2JzREGUpd
tXnkkHwfC19SlQDlhxTunYbPe1q8BGR1U36u02UGdsE+FbJAsD7R14T1TYLIef6h
gB7Y32RaoTboU8tQrVTXAJ9OS+8orpU4w+SJqJA0vpX4IvAJDeqOGGYWYht4Ueko
QTCv5bZEec1koH3XAqdyJ0ubRTjwOjKZvi4aEy/nV68HPQN683yacnBvtROljqtp
Eir/R/U112uNBuO2J71hT/aWEnziPUqEDxBxbmZ1s38385iI7tdx7mLMXeASWjN9
LGeqBOwTrc6i+CyyFFB6veRzrzgvCRrGQw6S4CZhaFKObwVl8nxGj5ciba5Cfgsp
4GjhbdtXN1Fv0pWuuxt0XjggocmroFnDkDaacrSHit+CEtByTUyv0CeUXbVyYBq7
HJ5i1FWOcdqlIbWuNma1Rd5hBntiCwsZncmNHnDobPKx4zxcOOm09JxBBIf8+k5D
uEifFzILIpliCAM5gg0uzBSLN5LKL6XRv6ZEenArePtg6AhQiZ5xRBuiN1RRR7oz
FGn2oi+d1IoD6WVeqQ5EYi3suT2+/16S/7077kVI5cfeEjxmb+5YlK32CarwJBHI
RefeZsttTwy56O+S2G4FhUrdycBmG7Kddp+3UIQ0TN5R4PgDCWvpUrwlFC8SPhuM
8rGRoG+ThinZ9qglNgZn+u7riNieTLtE7NZN4ciMh/4NtIu/zRoZgKIjxf8W/Fn9
oNE+5Hd6h0ZuHIo1y/xuawyjE2bNNmSqSveREYZ3Y7YkpiEBFkCjnAvR63mKes3Y
QtWGjG79U5s/FIURo3Hm310MvLCmrJRQePUO5bMDIKKwKOUAPdRIYtrt8DQSTglM
uUoWr6YkuCIVzwxpAD97lD2wdp9F0afkdAGkO4lEvjT9EK2yT8xEb76qCsuuNUQl
dWcIRfyjsrB+4JiXc0dY0BoSDvH6W5jn3VKRPGWnDCXbm37Utsm1kYz9LpYYESqr
uAPxdyJ1HmL6+k/ZpIZjjmYCSAhI8pYIteb6eT4BnF/edRdAd4WupSt/e6g9zp/f
Bm9ILq2mjNeEbIM2UYzbDnQJzlyPA5i0bRw9kfEtDLK656flHOVJuzqKRMrcByGa
Dop1W5V9Jaz8xOo3A8tAIZjCOG9jSCQL9rmO7jJeUBkf4vaXHq1Vj4mZIAd39m8k
4stYQkhQBTb7n49/bskdBBSbFvNOKNCVWU7cZou719ONH+G4bcnOsW3afaSSzOzh
x3lR3pXPSUHaLyniP03ncUAWP6WHKUZs8/BsEpBR/bZbe46QBRkAa3sDsyPZrZvD
ahNZgN274UFvw3uttzzqg0Y0nGQoUGRZoCHwTStckx7zQU+zZNkTYiYK8Y9zZPxn
AdYoTi1O3bNhUM/yMydBsMu40vJkrJwQi4DSOeasA6VkrBaWYaHA8hHyl89lKSUG
4vpHMuZziIAuB+s58zbq48WMwWw6RxI85gDXp5ycX+98bBXDlj7Hhdsg8wNBtmhY
vPhVOVlpxSK3l7hxvLl4S5qmSfHEZdKPKxMXgWBp8pT3howg9+HsviT/Nn0aB/eQ
z7GHB/28s4QV7AgXzTHMRRxX9cOMxdRB6sUewmatoESGPmLhKi0+arY61yDitW0i
HQkrtLKot/rHEEfAPuBE9f2qjgHdM8XuaX5leuE83EN0K/Nec3Mej2bmXtSSRsxu
7OHbf1eabslNOwvWxF8PaDrRfAx0s8QRoL2yBgms+ioFbFZPk2lDxoPoI4Vbx+/R
LRWp/ZZgxD2tmBqFrYmnxZwSixskKBO6QnXylx9ZoU9wYmHu3SR6tWRaJ0UdWIDL
yKu56g07HuuWDtXZ+8fzvD4qhH75QWGzL4S3LUr3DqNvYf6uwOPIKmeTHTVyHmcM
+XD2uwIwUIP+FvvA4u/6P8mWSMGVsanK2FGidaF417gmMgxyQ9ntPCKdkoISShbp
CiOSIxTxd2TBLz8FNYJd1tRylwLTfLM6/R4KD/jsTydDu5fBuvJLjLgv88iRqbhm
WWPLeD/KEkgcwzDCwisAJkn0Uijg60q5KGavNvcTm8I4vXKDjP5D66b4jX/cPQtz
N8QOO/kFqGWk4vUO2zyxp0O9oMHD8rYu07Y31C/Aok+GhjopmitegDTQzLG60TFm
iztw20OVgrv5tcBfgIn6wPznn3Hycu8D1RpytUzHcAwktJqNua0k82D+H9EeKxis
rzFyPUzlUfGpO87xanQqMWII568w+CGnQ1NmA5uPjTm1fhCQvZ+LPH12Shnv2pRf
BnGG/EVdmvehxXYin/c8ksuHYTJDZdTTywLRW89CZ/cd2ui+qs+lWLZGAfj8XZS6
0ele80XaXwUr4czq3691AYysV4rqhY9yUHu/IbKk0DwieVJEKOsw8v/71uIES+64
PSMEtNq0Z5ei3D3MGCbdqMnHJHA6pUPuMwWxy38OzXEBBf9OCEj77I/6eGIvvx/M
dcy6ewOlD0W8YMpUfAqvio9xUHbqcYvpk1GApEHiyoGq8+meeDATLIQcspicZOsn
79k6h0lIgU0W/d+bnvYQk4xZigNXEzp4QWEYO1i1AQhDYVFcsfg4ti/Nhq5GF1Tv
ODheL1Lbxqj6FqSj8n5sSVdw/HQ4OId4QwlUN+2wbA5ejC62bRG9XT25AGWXtiGq
qXrf9J8cU4saDR/8RHM+mu1h1uAiMD4bHoAfeUrG5pVD3kFYEcn6AxrrjiAX4vMv
yFEZZrPZw83MCnz4yRHHyK5mirAImeUpADuC4y4EZda2annXNDriI2MKEhJGNw3T
qErhkgZeguHFnfPS/Uznq2qK44EXwqsa/GEJ3gVvQJeYTfOPNGxLWw/L48Vuypy3
/ivsw0X2CmDOx7NN25/GjVHADSok2NJCH1dMUSLVDtEi92uo8z015dVyNEL02prR
tfNKGEEF39fgam0fyp8IHBGZSuYrdK184+iHMHiKbr5IF2ubmSvHgHyTnk2QUG7c
tgwEm6SP+f3WneFLmU9NwjSw2BG74JNLXznturgy5+JAe6Tj0IEX3bt4sskxoMs+
6OmdrYDQdFxbtIRpQzAk3O7ZDnTpQ2NTWBK/1pE3bPGP0XnW6SnXNRCnK0WUjGq/
7aisNsr4VLpXtRH32jwniTIaO5+KzXTQJOkliDiT998pAEdfmnCMx6Knb/vcGCbb
XC23yvsAobZk+O0goOyqQwTLtJYixRS13jjywnxi7U6I+ranVE2PfM7r7P3TOvYR
NzKWH/SqDjSwRYkTwnTjOlFG8UKE6LEcuAYomMSQIqo8Il/KqQoeGO+6TmbyR3fl
EWt7fsKXSLf/SHWuX/uHj2P3onjTok+F2P3exuMY35hcrmy4h7OnfR81oh1EB3bX
UQS9e8fQimy2Wa0lKF3tiFOjlM3bpVAHLtHMSZFVSnbrZJEtsER/D03rbd+MuSS0
qhSTwP2jcxep9fOK7q2igxJcuIxq95ACEyDdsXlGgMdS89wz1nstX57hUioVj6YR
1ZEaE8NEPhV2qUn1nQ0DRMDHqOFwicX7FYOLJ+eAZyK4LV5QpS9o/m6IW9JqqZLG
zuhJIGM1AXLTbphlVKkWGZ502Gx/5aCN8BVKED0oCse8doPdpR7twVvkUPDnt8sF
d9UJ8MAkznS32vkA5SnDqRSKj+2l9bSA7SA4cQpTZljxtrv0qGUX3ml6i962Hf+9
XkViXWWsjP7JNg3GaRpD8+6SvAHtB+iQWF8giTzWv1gaRYbq+QspOnD5T4BADYUF
xMG7ToqAQi2ivSdQyP+iLNYFgSHHfUnm6UTxprRyGmZ+mJfqT+oG7lKbHeqjl35M
HhdrNx+6dOnDj4IJVSMx14KQ66DksRmuJSeiTtf7VvH/dlMNgpiVhgnQjXEhKC1X
93RJtNugDxceNEmfKAcSdj1Lo24g3rrV720ry1DFmBWbe0voHfpJPXf1T4OKlp2T
DBqmQuxqbAsWj5lJ9KkQlM+HYh59y0O5XS2VPk0JPpb9hezM7J3GnAFoL+aDZf3f
j1CTGI5uVlePU6LXQEiPAWpeE456AwPqNUFMGhPwGAJdbZgWdyNXwninY2KXVcX8
AOX6ynwTTdO1zMOf0AqdIjk3rezG+fXz9lU8SaIwyvfIDy3ESuYopumVIpRjvOvg
BJaGQvUL7s89BRCQrWIkoWrdqTuDQlYfon0WnvQpSZnOtLgODZ70uhLmMeJr/4zJ
hAjWrN7208nOyUhfuHyrTwoRwa3gUW1Ud8s2tBV/VeUzUjOXgc4AtZvUKXyRMOSA
9Juz1Ota3W+H5SMV7c9Wp78VAwo0tJRAwM/3UEhokuoAFqS9frLbA5h9jN4brZ0h
u6PXeHz6I3PfdNpDdeFZVdMEuYOtdAlzPKoOYwM4JtVsDtj6OiptgDMhwlwtzOlh
+48T23KxtNr78fc6r+WupKY5q8iSO9On/Keisowcoi3LQwoHNojhh9e8Mttn/ahX
J9BiHel6++DdsZ3j3RRs1ZbY2pOsnsjGJQ1AP0OKmWXS0OD6GlWc83lk1IA1yW9m
GC0UX8OT+BuWkI0SGH6dXw/qJHcizDViDWu2T+gnkWa48ugUlRqAMw4Zb14tWzH8
cEauDzdrqBLYIV4K8WDet84KiOAJU1vw13b+6RyaKrSCRKnD/VhMQB81RZSZZCxr
2nbhNilTMZTF24NMjV0j2+JBpE8aLSiWlA89kL0BwOtyqe6UAaxgSq9/A5W0C9p0
8ouD2biufgJrM87njz3ZlEwX5Yx2uVByfg+vmNrIyP/Fyff26dGakLhqVJ3i2c3a
qqAyg7SAgvlaS7FyhLqlcS4mQD/P5ers47xkJSGJ5PbFyDxIchUhyz6GcXBDVsMF
G1A/hrL+Hybrzb/q8UtjT8wav95YuHCJVj6Mp0z2ko2ZbOjIG3bDUk6E3oqGKpku
4gjhhujl/fQoAue1xB6zjq9ucI7aSB5ZNb3KzRdzyg40IXMvVHo6hZVdGXrFkedz
f0h9MPmy5LeWhiSGHVqf+cHza/drTi0ZTy7f7Oipz0kjoFr3VvvqJN3UupJdNOm+
l3725GjsS58HAefrkRxxluX4/e2hTQL4S5mbeEs1khJrePZdShtbg4dFooeqrOqg
L8ev9gwxNp5EF1gBgQhQj7G28YcsagIWArhiXKZnYDARWuYVgDciTeFCOPc3Z/a3
8dI42DiG35a7iamrvX9M4EJz+9UbbQU10KraEDLEka2S2p197VUqX0GR02ipzEOD
S+WtREBx1isVUSIiyywXoAIfMwBIwFQBJc2hAU3SoDSpOQRYcCb5hFR+Pym72s9V
qn+xE8yWmXwTq/nYbwja3kQJmG22XlnikATmttOTUmvpP4J6BeK2e4XIAeTVdGk9
LphKcxHI0/Q7/rMt5BwN0baY8ovwQA9W7kMbiJbkHRdEZV4SLZZPkMNCkaHoHoQw
nnIAXwe8uH6FFWmVoan4kjxz6+GN+Owaci2GDG/n9FZl8YDKNAVopI5MxUid4zCZ
4KM0Ya18ghvDNtVKVnUZSc6mKxtrIHHz7w0+YA1FWAEtIbxfjM2bk6yY9k6MPxvp
fbT/PaZJ4qBtIVF7fQ9P+rkVJUitb65IMsh+oeTrw+XDFyPwLlkBW9hVMWYeghll
6wPCafMCUrq2k3zS/AToxoKQFhmN6PcB6upzQ+0llM3CS+iHV12PUrHt7mJeG3QX
ztv/UjniZ2xfYLJImd4nMrmdcJmamAscn+Nn3IWhI4C33DsYk/yuyRI/mBIsGfFh
VEdBW44qaS5ot6zKmb3HoySczDmQ1VB48T7dvTKQ3Y1okEKeujFVsrrW6LIAKFL5
Y+AGO9mHEB0LGMUIgc6eK58OBf2A5NeOkN9mi51Z4sHpHcRNreVQbMQfApy4YPSW
e2MZniqrS3ivHHRgTvfiQ8qD0kO/miqDR3Tu6cUlEBgQcB1c/cPz5F19OHuXbrDV
j5ZHJdgiDi/xU42zJXxi/GASCCiTvigbf/9vRUHAzPx3gyTPg0Qg1XAztflFzj++
eGaHiTV6Nhe+00/SjFWNQXmCvFUJ+SOIbPUbwrcTGJ3W7dyF4ERx6swf0vsYlF8k
vuinLz9MlMB9mZ6sYKbDsgYNnXuDP3XFq687494ss9Fbfyw3vxPmwsE9indIjp3y
V7oUwzptPwYHt7Gm/2XSiroZYQDZcu+QCyN7NdUaLYNrU/lseiG5V8qq2Q4nev6W
OX1i8VFrwqYPOdVI/adHO78T2peJWcZobfN96dBcHKruAn0S4OBCIXMYvhAtbzjN
GTVrGFznaI8ebL4yIpDEA3WrDILfFty2IVdY+YWHcSaieBQNWrQoBiYa9/Ku8fhe
4pXfTBBaKxGo8RHGBgUXTdi/uq2Wb/T7E0sOK8aEoY+smsPj+aS7gbGxkY/uOyTE
pABnzkiLwLuCfFXwEN6gjeUpTxRolOw+uRB27ViVvGG35TwXKovGVKu0QytE7usT
8UMMyGpNn7jcZZ1n62A9QyNT2iatU96/yzX3oog/V2yn08AI/+r7pb2GEy3XZxQv
tbyEIjCoHh+Z9DRlyzuC5n7sFePkpV78ZzFZfLw/wNNZ+qtFl00YmTq5JzN3OECp
Drj4leggUIjIuFKzhuas4E5zot9EfSevMoaVlB7DnY1D9Uxoa/73BjE1eB/P2PN3
MNf8MdlbdX9wq1V6o4uAMUBQjrZj1Vtiaz3yt1dQ46NLP8BJQtCUZilEFlcIjPlg
EjlqDMuklWjqCcWHvfo0eC8eEP+ssDdQRNgt7vvJhgqi+RpfkZO2vN75qglGRVDh
Wv+o27iyPNhBBGPu46482kjUxs2gGuUMHZUl/dndssKE6FyPu/MUTqMUxWXDByp4
Kzi5Ufn29NXFvVrZ2GIRwgv8mQCVtzRYP4oU8kidt4WoSJkyI/gEvSGO0sMu2Qem
HflFtkcKWRZjaDFyo/a22FO1+dtTBJciyC7b/RoSNfzkAxht9LsDn3eu8l/Apyzj
6cqt5ruaiWaZx+k+uGWN5pkvR7KmUbCxR4YBsf2VzoDXVvYJ4W2eYcRtx+UFLIcA
T8xtjpNy+2j6fz4WNBBJ5TfG/7+/yulq2WovHTa5IYym+mEiZRyUDqZzAk8gfF4G
T1C+H3dSDw6mLNInmFn1ldG4EP6/iZWh+oVlAG/R3mLH0jx3FLgTIJRaAm49Jt08
+ZDu5FV7sVTFxVNZq4dqK6f3QkdTxC40eQeCtsl7lTm6mqdjQUPDV3yNsCKWSR5y
c923D9IMG58vMwPpBF+LesIhS69O3Aa5UM7fs0ywvB9Z02yTdgkuWTs1xIQ3W6Ty
pLvpx49wHdk3NQlQSeYZPD8q9DO3KEp2mijsq3HtOsGR0qpsl6+189UWG9C33gwD
mgm8Gdgr+aZKlgb2Mow8V1219ec5Ppyp7QKRWSbWvmleIDkswrdbMfwpRNZmyE5r
W4CfeeUB5Hv90z8P4kttSJc+Zir/gifF9X2r0rlvtlFCh4ShC7yPbuwz2bFWqs/V
HzeeYvtbgJTHBW16T3Y2toVs/TM1fxYGabfxT24MRpM=
//pragma protect end_data_block
//pragma protect digest_block
YnPyLArYIu1z/6bpsu6R6So/7so=
//pragma protect end_digest_block
//pragma protect end_protected

endmodule
