//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
jueJ3uGbvT/wIuzp+SPctxKFLdt9eWKFRHDV1OqemFFBftHXBssBuN3nAQhLm33W
EQnLkT2WyOJhvIeo9LPi8ZY/aFbZO7sG6nJJ7sEPVQS6GQ2FrmO7iuGrsZnzOGMZ
FueryWWwAD01DGvX6y2TB0Q97h0B+//wEsOAeTEz8h8+GXN6EypitoAJj48l6gjv
V6Bwoo19voPK8tXgIeUn9Nkir/2RnOF+YyfWfT3JX1KCcC4jIEWM+IPmyoTA5Cwc
45RZrnipHW0kqYi2gDHq8335pb2s3ZDpuQhGHpvetuWgPvWPKNiDGtoivD6cOKd7
cb6lfFkmxEH0WI4y2lWdSQ==
//pragma protect end_key_block
//pragma protect digest_block
It8iyQP9yfqfd+SG+Z5Vv99NkOQ=
//pragma protect end_digest_block
//pragma protect data_block
VwllPnXcxbxK953kNtrMqIn+YoaUfZFcoDMr2SfQ5vVWtpbYfHH3cwOovaossK1w
Wh55NauFpswSz2MjIfuEdn5YEQpb8dg7pKZYoXedkkHfKBhRZVzc92HBVnAYd94t
7d6tx5ExrAY3gJundGozR2Rs51jl399NdUxZSX5KZksGG5GyDW4wnaNmXDJcSybq
4xOVfGUZ3WF6tT1Ay917NN+9G10k/Aa8NhcVK2nJdpeN9aIbWzujfTHdRZC3zYjH
HtYA9RdQyvigyGYp1LSi2EwpK1RbU0D12X/g0297oUEDFrKZlEKJArZ/asssyTsk
p1MWHxgFp3u0QQiA0vNqnPU31d6JPr7cfHdNjF/oquNnYicibr8MkMi7TrvX/Z31
ZQk8WYgxCbtn050dwdLyqi57oYdvHzUuqU6Ljv8xvZH0DRNokM+t+ZGH3n2zncGr
//pragma protect end_data_block
//pragma protect digest_block
ZDaQqFsJa2Swbbp1wWmSqNrXozU=
//pragma protect end_digest_block
//pragma protect end_protected
	`include "PIPE.sv"  
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
o8Koo1LY/A2Ebi5vZyB0T1jy51mnYoXdEfLRp+S+CGqvanWhhYjNOUyp9U2sfanZ
X4jBjxQZY8vnFiNIIKd/oyUnd6HPOPZIa4pcWOrPIQsvq6V2puXWiUJs75YNaF1O
li3g7yCqeGZpyoAOecfns0YjRtCvHPZwtJrZOQiG72PtVYoEYrNobVbGAihLoQUM
AelEyoDdM1yyfmtNU6SFi49MVkZ3up81X/FluGTvJDujS9VPTbWQmaWdrKY0acZZ
y+IgZmMAcOoCszjc+mLHVASXyO+F7d5ZWGxytArcNC2R3v2kSc/0Kv2rofwselTp
JBKpZNHhYiCvJ/+6PM1VFw==
//pragma protect end_key_block
//pragma protect digest_block
Fs2GN0pXPp8bHm0nAToJT2iHbl0=
//pragma protect end_digest_block
//pragma protect data_block
kWHS8a+6dwSlGEz6ykfFXSX3gcAoXgyTA9z84AXZQDolWYRpZT97iVMNVPtDIiik
W4VCuOT/W0a+HrroDUjIKGUk08X5BQmqNdn6nzkZjd8UNGNU8v2l7seKN3QIs0BT
2Jz9Bs9ZeE3YGpB/QBrc56Eqfq+iDVaSMbhyigfNNhjujNMqeRPqfk2unS7Uaa7d
fO+lJSeWlA9OHSH6JACE5He+2mihGgN/vPJrj/YWe85c81CGTsmmKE27YUjfm1q7
ahiWZix2zohO0sNVynPOcjEBPYpo4ZuokrEo3jvlrxa8UtrvYt2c9O4WFkfKWHdO
/Uc4cNt41xLeSsTOyPTWz/GTAqSB8uLsDycDdUphE62qSXbGUVNOkHO1OsT6Rf45
deGf1nuta6g6nD9w32nvN28JB5kS3cKFTaFCwL5FcKg=
//pragma protect end_data_block
//pragma protect digest_block
KE20oWpN0gkig4M/NzSaS9ny51E=
//pragma protect end_digest_block
//pragma protect end_protected
	`include "PIPE_SYN.v"
//pragma protect begin_protected
//pragma protect encrypt_agent="NCPROTECT"
//pragma protect encrypt_agent_info="Encrypted using API"
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=prv(CDS_RSA_KEY_VER_1)
//pragma protect key_method=RSA
//pragma protect key_block
bDEFDJjBMdDGHNZ+JgmU2/9MCh8+bCaWSt0EMyz8oSKKrw0HuRn4Fx1Ihs00YlMT
alKLLJIcDz3T1bG2S2J1VvduHchN0iLMDVfHm5ZWBs1g7CFHwH9aW++1RgjQsEb3
6f5ym+dH/xUfEEK94oXMPP2/Qf0NiSWSzqKa1Fnk5Jt/5VBmWzPrptoOST5qC/Lv
lGYnXQhmS5Nith5T4D4MOwBQPXyVV9r4pOh0JMxfs1Yxml+rCKIveqhUCccFADfY
cAcTmLnRJpk0+0HwogdNS3Q4guhwDci1Svb3Dl7tESKjMdVZNBYCdIVic+Tg4abu
2dCXM5kIJ1rkleO5g40MyQ==
//pragma protect end_key_block
//pragma protect digest_block
1NFMDK4IRvwgTKkwa2U3rA1tluE=
//pragma protect end_digest_block
//pragma protect data_block
lDwHuTc9krS5nMULfQto7NXgevbQpNXEx+Vwi+2ZEMCxGbo72baCgqrXEjKyDHcF
TSUYbXczc3mC/fk39FMzn83kCAxFkvYh3dyR7ghr0MfFg1EyrTZABctMlJDHKF1O
+hhhmBxPU3iSO3PhUHpqum5M38+VqTemeTak4Xxsy8LSxgAa+RofEqeTPR3Z5dvN
NJaiSmHTNIY2a+ioAMJVfzXJBoxAsG9Xr8K0ydkp5XpF5g67V/k0dZTF3IbZTjKU
s0oLt+eQSfLpLWg7MEQmUH7NXck1B/pUwENNBmONmKXPFsEEs/X3L5Oi/wgSVois
RVR8fZV5Z3NddBVPGQt3WrjSHyB090mk5ekb6A1dGSKHvQ91X26kZooSTc05kgmQ
Zozt1MKf1SOjJKlQfQNOKfrToKMb6Zzw6sX60nO0VcrsiG3d8xt4tY5f4d36JR+B
JFxsIaZCdBoDZrDNAbT+S1b3DY9VHlw6cZs7jmWRM2nih341mOq4EnV6zqlcXbxQ
1yf3YcpskirNWs3r/HF/xwqF/5GKocHdZtGJqjbSQO+Vwd+NSJuadLJow4BnLCS8
1onyaZf+l9VPXbxnHC5N0B5flrwPJtsMIzjWGZit3BQXvDnX5B4w/BR1EWY034J/
ZA1PfFEGBjufXDImM1vR0EyQJnSEkn17BUcRinyhJgKWh8/mlWBqP7o6GNcN68+S
j8tE3lbcwN81a+ZTrVY4jVe6KNUWCy5mxgCy2ihrvy6nLjJwZ5GngEc9PrzUfMmZ
2cbGZzuQEXM7J5EUTbbH405Qnf4jPVdLhiLOPE/gy92emgvWYIM1KXbgLldiHYwZ
rhcz7J0pkZ6XTShpRVOZbLZwd7SvW5C5B5f/zkXs1PueKUuCfBIZk6yndxfFPGAm
5pCtMP8EX8w5uNqUc9df3Bw4EQTmw8A9PYVZYch7AQhhqgJa2gjhgJe77HJp5Lmm
6DNJxNV24krnQSmUWrNy/7Y/NKyEN7Ne6iTNRR/8jl/7Q9wwvwsCB0ALeEeJeOnF
5ki68N9al4JyJ6UKo9igASJczms2AQ/5uHZ9AlxO/ChNccQwXE2z9DDImPVkNJkE
AKD1906h+HTvkIoEV6rKlzrIxeJ+SvBRCR7NZOMjaa7PyOvudxUricHBbr4coL5U
ZTYyL4Qq+QI2jHwltJ3xRbpqTFinPpkNUMVLY7I9YZOpvFs6iOgfKy2Mhd5qehXV
qQlmKLLxXK6aHpfBmDIrpcDrcZdOB82IITt62yb8MxJUtaRydHFMteMv1pqnxN+i
fk2ZfHSTHrmFhKDk3TXz8WX5X11wDPNt/1/Xa5jY/iJk7/Az95gyX5G7+7QotIoi
EkaC4oC0+g3hoJzDanhEBccRohRhgEiFGyymV9hh2yZBFqBf3eRqvbHFBuIM2zOT
Wrl61m5k1VQt6s8//D+rqk3kBF5GP/9+bIcFgbreZRvKRVYjmoCJjINGqFchyF81
AFua6ymqGWMqU1LVs3mLEecAUEJfE37eTSXNe4HiStqfY33g9wKA0bXfTfFeRzyz
K82/7VIeRynvqAPm7Wu65PxcSH/++n81FBnrve9RQRauPudtOE+ERMREZsQYhTLr
3pGag/KoPnC/ZAtIUiNf2qVB05f6B4GAyB7/N5u8SCWfY9oD2fJ95Ufrpn+ePPZi
MG3evmHkPvLGR3Bh9rqqMq/l6YxHypSNeykJmRjXwNhvXF3j5o0wNMk2maF+9UJU
jgVxnw7RpP+prCKmbiBKcYc3lHpEsC/79wWCDMhb1RQWQ5ICqRMPwJ2V0owSExEj
KGKrOAkMhZv4j6MrsdouTgutNZ5KT5+Sn8HqAG8klDDZECEchI7YuP1wmcEA7XXO
roUH8dQ6F3DJZ7ArKc3QZD1WVRRKInZ7aAfc80IisjUfXtUA4gJZS4t3tGk6oRgU
cqDr5n79yMZ4j/OlcKXwU/VAhn2A/Fx5vuyYH/JwOcpi+K6OQghXEPf4WWsuZ/5V
xoL8WpfSkaxq43a9teXwU6oqC+oz1xeT8u9yCbZ0hvvxhwIaiCJy4YpqD72P/gk9
bQIuIfklGH2YBC6xnijAt9kp6fL1vDz3DrBTtPpEZWIpfnV1Iy5pfkyDBKYeQH+E
P6Pt2IFUMIagkaKlIbsnd9EbuhpYnL2zw8JzDUlxCrJ4YhYGEjqD4R9XcpLhXS3a
EGKeea9s0VQ5lZjMcF71aW6cezWxhRzfxK2ovQuNO9ddnxBPWxtEHWFl5KsuWVip
dPVlW3vQ6Sr4+iS3rgtcLpnN0d+HCdYwqV2g1Pbjb2lUW7C48Rf8wdqu4RnxtHqO
VPUr9Fdna4jvS0Gx4tr04z2EgAVWAvtDrlOVaE8fb9VeZBb1gatrQULAc/OXyCP6
TzBaTLbuI5V1E3z1Zx1kSy8jSbPewY26pojUzmigEn2Echmm0F8IkddKFKd7LEKc
hH/MSqF7cR/ANJgVru4qJFEv132hiO/Qk1U2QugEqK5tPJSfg430JYLK2r34NdnF
qNaqSRLEcm7A4W+B7loi1mvME9E6wMZF0rEsxIo0pm8UgCo9NKm55pc5ne9jS7fz
9nq7hi7EOrn+6EQk+rzFSYP7EV8Te95Z3IgvTZxcQ7btZs8Fl02he625BLKtdYlu
zsaMGDGzKqwth97ZWv7v0LHqHcrbi84JVdX2LR5MY9P9dzQrl9vMxbzb/tZWeZ9t
92kPyv2rAxqcpQx3JZRj9JOSToTcUj2dgbXwbFQrDUQx/bOryt5jZvWWLCfRi/AF
oSu8Fjb6n9Ve1idNvI8TsJxR6rBC7IfbvZXo7I2AIDnpbabDeodjCEK1nhhVHi/A
LSJm+lMfd3DSP3Y7zRGBNpClM9GZoPs0Q3Y40cxcamC6c2EN9IELgYxskZ5SUCce
mmBeBZ8VagFTSvlyFiScgySqHIQT6lkyIqfcqjPVAW7sbmYG45uXXIJytRiS87nH
SCQlluw4Q47pTeR6wprZowd222Tdkx15LVsFPiX2ZUMIPcFBCewf3y9CEIZr/z9U
B6fmkXxOQrSa0UrW8vd3moMXChGTu7FjNGN8E1Iayh8wZjR/M/jW3pndDVh6wzrG
UFRDrj01BUQYbrmSVYNUFG1T7pizMbTZMYvxGU9GjW0c7wbBk9nK5e7mIbVaSlgh
LEhTjeWa17vOX0NjRvqnYlZYv3xWwouHTzBqeyo5uj2pX91/SIo7Yl3LXE+6nse5
TqvXpKCDmuXsQ/qXYsc/e9+NknvpRf9nPl4iSvAIol/dToRvyG0JpJckjrXnygn7
rT+3/qrvu+ZiZUOgc7NIx2REpR3Awnmqu14eNTxvqz0s5Lhys0sJTZvBlHbnZai+
iWhvXGPcGDzHw4K/Q0dWfjbyWDId4cTsidN1AMkHK0wo5/XlN7aVjw4vLssa4ZTu
8hpIcNz+k9GvZfnduwcvmTxCkeVThwR/nApU1wTdEhFiHpIOWpB+kt0NTAwwETuB
6A/4r/RW+LF4jgfH/PjAP8R1cd1tbraR2mMG7HVTKKisUGWYmlMrT1MEL7Jzs2Z5
t8TV3/VYPHZx+dxezcTqJeobrxrekFGzPVVbwcg9V34pJ2G7HfOuPsRdA/kppHdN
s2pI7Wxvk6QYUJteKZMH2fX11BvHWtyjoAlrliqW02U9Ywqxqv14WKACVF4SBCS7
Bs9vKXXwdHXeZFYPICFe09E1mJQvD7b6tVUHaEG9D3vDHHqZQOzbqHS3l/4GToHh
48UUc2IB3nYPHK7tntNOEtJd4iFud5Ua4bsZ810cahyWzJOl3by2z8nF3je7PpU6
SmEwvajOIJL1qsIR6l4JI633eVq40QDL/FUKED/laHaO0D778TOnZMqY9vw70Cpl
h4xbB24HXLGQyq5RjvcYHvRtpQT7o9sVrnLr3N/my1N1HWTQoDcRxdBv0y1labg1
xPjD/wfwZaXhEZ1y4augFLZ1pbqh8PuL3QIr3tdss7yIKxE7MvcQfPzgFq2kn1+T
yvbw+4cJRVs4E2mdfqil1iEySNqwq1TlWlPfIqidxqEm5nCWgdaTl+SYKQGZPAeN
pZe1RmY1HjmGlEIGPks4SMGwAwtLkWrs8KqXxyOFcOanKA8vBflQGiQMoi7jUOa1
5uJA4Rk7Ryw6IVdqXITzUK6b9mQcHc+C6NBgbtmBsS6ladDpH4HeJ0aX9DrP8k1S
CInNnZJrYN0lcqPdUhjevJTn0ld4xjPiZX7Ad+Oi3GvDqjY3GpvONq7o2r7hekqg
kXMy+CecnFnjz8Vq4pSYFkl8ePT2kBf1lVjWt25jYrhDX2hAz1SJckBXgDm6zCBZ
J/Ie2CRCAv043AfZTGY7cOhuwuXYUk+lqSJEE7gbH92u13yVdCagVSWOU/G9pmjW
KgKX/sLZTvcJPYTajgxK/6RnIVPGEJ/d+yv67bkG8SZOFQhqASsbbEaNtt+29aA+
P5roaFTHZ0c0fSgbxpFIfcKqzV37lo76AWUUOOVq0IM7UTAGMd9dUqtbO52Hm19s
6VmtBW/VM7yO2y62K6PCbU6zPNlTpO4wqPM9xQzpCCP4JvB6HUfUjQaQjFCcWNgx
5mkSD8hOM8teY3CtAy9+1MiTW59H7A3Wyt2xuB4dixgFUvVQJOgZZyFf7mQ70uTF
cjQ5RrJ58Jvcl/aPvw1uRrGCMH1LJR9+RN8yJerGEr9CM7SUm6ri4U3Gi6Nz8T5o
GtyqnVMvrO8xhBAi2Y8B5pWzqH9LoliNXyhh5o5BDth+mVawJt2PIRLd6OHPtEkO
MSkA3t4AjR15q/7f9qM4qcsEu5Zqp/287x8sONLhAbrvIorY+rqvjQdHVtaiYBV3
r0+4iVC+mwKWycNcwFoyDSVlJM6hFSwnFf8GksO+2282trGvuT0uQBlh6cBSnugX
+eSyxekZIYwv6QrK8cKXZBi3lxd6LXal+4aD4IyHP2NfuizqMFcFLIdEON0TxNKm
itpfWmMfyyRFbZ/jnFnBq2XPLCrkHp2WqyWZBdAulyPOA5/EZpl7sbYKE4NlEuSe
dG3wk2dSteJsilgA0JV3EKyl1KO+knZ2besx2oHdpgETCpkHmvbGwT798UUwKymx
AFRmvai0MZPrEfExVtZgdUIZLIALGtDxJOIRk9ghsug8EDUYVcmgKlR/P5e2guhF
7g/PZtsNGNFHM2inw2TglXr5/fhkP/niOECYmo224ecLWjmrdiKSIrg4JD42Z8gJ
yrgQzaSJWU0++RVhGEyo+650vnIzqQ5oGeztcAGMllSfn7QYre0g4sWV4Lf9HCeI
veN9sm/ihcvXaDMlIgnR8QfLJYYCC63XyvxahNQHkq+AwIjfhQ0fdiaouWDk98NX
Bv53dxN88J+3WxFE/Bu22CfY9S8Z9joyWTJJl86teXZWrayzIi7fGIlw/E4lUeJV
rtGJBByzTMMBwaU0F5IjAVLFmwMRGfjuXOLJL61K3wN4v6+vdJnaWh6iNKAOz1nh
bpTlho1F/GX5K09X6sDIFLUrdoGRxfbcRLN2hbjy3YjPFcWXdLzwr1OgJT+jcESE
LgRHcwQIVKgj5VVQ+/CGyu9Ol9pHmeNzkaj+rx+G1O4qUUQ97ThVd9HMwpd3EcK5
5/ADEDoIft1eW2tx1jfyfQAgkeiGJa/zkc29aulaz9PdH692JNS0YhHmSUAz9n1x
YohM+gXvKY2Ljk5/GjaY2rV6S2gsb2t9Rz3zacq8JbqiA5JFxhxt3J5kYmQ1Iksc
TNPP2stEx8oTAYQ5rkZ0oss0IuTKYaE37XZ657GN4i7gXt7WQAH6tMhChcztZQqy
0QvrTr3g+6KDBAkiSVNlGR0m3OQdioKT4DHnKpZdo8hWrTNI4LLj6rV2M31YzAaW
miDEQ/n/jM6hm2txdTFjQvDwhqpph8130a42bXhB+5Zj4apgV6osfBGevNiVzgH8
qs2WQUbm50Ue7UJiM9YED2NITm4FQTvNwn0IQjYYOw+/JVkvXrWi11EccZU/kVWc
WIe37wTsUk8UjVVqkdtFdetgukwIF5oXJ2WRHcVysuxz1C4n6WtaxXT7PPpWCSJu
Vly2bElKV94WUT7FQo1TXtW+Ttpt71muFTURFKcjottBwKba/EegtolKHqRLUpGT
6zQ+qysOJUxLYgSY1GLmAT+hP32VDWneTB7TC1mpMqBsLRARPprqcmg8O3IYzWJT
vm7oVMcHASIIJ98iYDAgBHKoKXP0Lidsm675HaPquzK8gJyvbl2N+lyWPQ6z2YBT
AjToMJcOi3baTwHhrxLGj0kdjBrMKF6OnftcCtwGEixvvp2Q9OuSgpp/uema+w7T
njto+BLUoltYmrFiNnnA5Gw0eB2gAOZiisEA66ROIWodvUFTVo7Reds4uIt3WuaT
tMd17Q/F91hRWyVqv5bK8y2tMX2ZnPcQLtQkc0MtcwWmrWu/ij+CuX+B22UxsuPb
UYjIc11pAZnnE20L1PWZ/THPDvWxdpA9Eg2nDjUzokrdVShy3q+PhW9yJI8HnShm
nVyHcVN9bmwMwOnzEx+0zv8KOl86gDPF3qR/CLhgikU+6ispvBSrXOfaqyiwaAvW
/CLu96LHNBghipD5x0g2TL9eGG0zDqb7XhqJTJ7EKvEE/Q0hhuABtYe9q72D4f5e
TfwtkuXKpIrBimhLgRP5xBAorsXsU7y7Jiior6ZksU+35RsEhWQobohpGb5YB5CS
8EH6okQxnX9BXVXa1PTkjaVi+biD+05JVnbsBnnJfCQfSS3hp+0LZTYOTT4dsO7H
vMsd9hRwjWAqLnk4cGcKQlw9cRogMSXnZbc58xEsx+EaY4/dN+HDfq+S2F9fMomr
lea6gJJ3zpn3DSomh1MnXBzqGLikK/vfpT4ygunTXpFSefoD1tyaeMF6ZJO9hyND
wFuqTHhVmK2Il6RE6oPQuC4crJSqkmpQYGdS0lxvNZ9n2CYjLBlgU+bTNFA47AXD
damMVfxPhkDEdAc16qXNCaxXSfhH/moNxzzm46gWSlEJOiDr4wxU+UWMMTFBxm13
ipoI5SevXZUItGFIdBm19+3WPqduWbDVaKa9g1SnTGPTYosi15WjqyAkFMd3WVaU
It4CTP4zGDvIB14mhSoBJ+4QFULsa7Z2qFPN+ibTDdH4aIzoJ6kGpm8LWqyjbg1O
5cLpuSCBtudvQBL35EM25bmhXV4YLcBeewaqQHffZGbwLhUAz84YA++rOy88dIz/
sXMOqNvXSpVvz0tdmyFcgAMs2D3oa8TyAoH0WL8aU5KVVv4XQLhXOngad52+/57m
YCPdqwKIKwOpRLTn1hbluUif7RmL1BqcC2YXEjUONVAoEni5ebC6eRFM3YJvWO6n
Hcw0ibk5VNMtl1pRVON7eTzoXVb3bRNQH/4jVYNqQ8j/11vjc5JL1sm/g8kHEixd
QAkHsaXUYoPB7/ZBCAtzeMhkwV/1ncFlGfd9yyKns5TroDXW3pvYS7MvWwnE9J0t
b3b+9viAcDvMcwAdvGrK+r++AcfjSWZbuTj+b8wBOx4qFVe1TPEzO/RUilW7174k
JpzryihENs1wBXEwuPgD8rnib7htV8BGxlQghLJ59U/ATP5yhN1wmko90bcPTfCk
uXs48duaLjQAsGFdBJ7dnyhzl3jdsZ5d4X8AjUAQBkbukCTGbdnxw3h0+tBx0H62
zw3Te4tONinI7aA5BbmDG3XT4zPGFk6q65ZxCosEWcR/r1zMSOaiFoy8cVAY2JSV
uyUpumtenI57SBjs3BBe2x2Bt/in5CQWM83BxaR49vt8qYh7gJEXOyCZNhmSVAKL
Zdpk3kT9KCQMFEJA2AFHRv9ZDLMkzvuMfTl/NNs+a2TvO2CcevdowwUjocKRSzPs
hdixLjtTJrCgegVfUz7aa5u3x0E/u3fXvQxur/o5YDRbrl1TYPDR3RiYNDY/S+vF
Y7OEVbZmPw6HN9c5TetrvDzGbhYKxs00sKZU4y3TEcGcsQgetYYdEso/VgCez3a1
/ONoUz5xKxcLji1qcsiYCkq9rt5U6YToII6wjlC6S3tMzEkKrw+OWB1G6ZT2LPO8
fanzjpp8jao1DZYVTYcrqs4d2eXycddmSJmjwbsgyEkOENOp6Nn95xnSD6gmW9fP
zhH1Rj7l7d+ZfsNRd0nhczOSDAFkA2m7Vsz1QAHURGje5YuyrZri9lM+PhFuML+4
2rytWs7FaB2eZkdpZskVGHyWpqPyB0YjD3poOqWg1sWbyMCBCKRStmaaUoyWYk/0
X32TAEcCeTcoHV1qlgpYJXctloYrwAa0t5BoLTpPPi4DV9I8EsnH7gVzLb1t67R0
THx83g4YV7G0jh2alL5XUZOXCLlEPzjXSROHth1xWQVGbrq4UqlK8fGXEesh3N3g
83Kz4UOdEDw/OvgGMy7IQnClb/HOHUZ8DrXcOWFRYX9OP5zaRmb1TnT+sjqFb8qW
spSs3qc9C7pZNUWOVAY9UUWGowFoPh4VpbV/6Dr0C+wR4jcwn9AvpoxUC1kfrqFD
6L//grwi2yguOhawRleTPJCHl7m2hqFtJIJ9tnXGYZe6jI2z3uBkR4gjmztI38lI
/K5OJSiZpwXd5f6rGNAQ90ZjbhsexpyDMPSpj0SsgiZkrgOyufHZ0tBUIO2K3Zok
5Lftt+QFtyGDRLvYprX//JLcNzr6wIpF79a+fZ2zn/3ZW4P7Mk93lwPNg9+ptyRS
fqRhWEKa6R5oHMv+xd4HIVbySQsj/als6e6K4YY6Xu2Ok6nOuYWM/Mot0/P1Vxl8
aANjRsOfEyISfNJ23DDPwsl1Je8ps/BBNDPjAuECiCS0O+xvxY+o/G0eSehoMAiJ
ejRRKcaNpoJnVEXQfM6qtbP4xVwRmy7hulSUkfeU3jC35o0R5foSEUwIz47oq5Sn
uomdaW+HigvVKuL0mWu8BFX1Q0uUbxmbPASunp2ECcgMsmBKvdYozOpK+wQWIh1N
8qygd9G+IuO/RkD6le0PpoQzZSnxN1zebXOPHc4mPh6nm2LnOz8BpK9pFRNAv6kP
qwxGFkIqzlbIMnoHlA8nGOBRRAL5na0QlUYE0zH374ZGxTWMR9lbo1sBoCWyRN9T
sjxdbRHe83QYk8DHmMjT7mYbADuHSAzmSbodpu0G1oK87ZDKxdUjL0+MBl5WR43G
406eGo8Azb9RtCKQ5oZoxLI6BPJmHlccehu73Co4RWF+Efjka4+7/lotIEghQJ/y
5p7q0UQ/iRc8g6M5FvFji8a41cujI/Gf1ZA9oyhVIVjw6O7nTjecJXtSLVwHj4Ag
3oB5IQK/fx8f2nLbs9gw8EDNRL5J7yqqVnddH2HOi//RHeeayhgGAampTcS7x9cW
Eov722pNLZtUP4pJY7KTfmEwDsOCOWcFCd4rqNz7/sXjP1q0BraXPhM/IRXY3Kgw
TWosidWu58+dTM2fwAs1LUMfWrzEdOVX1OJ4UOgibLRMTZdAm4OD8ILmoIyRQFZ2
M2r3J+XKGRWmwwGRgCh7XapYqG8oCERM7vVTBGwq5WzlqmFSUeP2Y47/DePHwA0h
wxfpgrnhPl+HyefYZeL/tm0jTasgddkCZScRhJqzq91HvpE0egZlbs7TB74wAnPA
5J7xeUftSQ9eQdITw23XCk1+W4jvWkDaE9t/RSTjPQytBDhoh80DXuoPOaNSsrR/
X6g0oy9VzOl3tf9bw6s8xbiUUspjbnCsrmZLktNHvwg5paOiphwVNxFliQswrLHF
lkwU2SV160+KlTdjgrm6u7MjZuYJgP+SFLanoAzlqj9g3nVa3y8e8eBpReUdNsLU
rALpJmLfpfyFVij/bgImgtxMK/VhMyV1erKcJWmSaC3KC9x5a2ZxdB8476vjgXxn
BQVFXULHYulyEPSuMxDKzqBUiYM/AkLSEWdrw4c/TpzAyiVYmnAjAtW5g/cctxv/
CzyggjhwbNOySd0PDDdmsgC59JrAKqrRsGZjCGZdbVu+WZaD+43kYGWCy0pQ0Mbz
ubka7OvZRQx21Y0H8jNjlqRoQODqg8rEHimt1/H/whY/lnxM48DqHQIH6NSCv5RV
7cGDpFjQUP/ij2YN9el3i5P6D3gfE8+oJ3Ls2pY22g6U+GYp/y28kJio6jnyQ/6r
fekzO6KeDcBJ1wxJmi237TnOfQrxOWMJlywB96NmNmd0rEKfs/DU2qJpk+NWyD7M
bMsWvNZAuekDlCqc++B5tdwrhwWRG4UKQwUHjtnspP3R7xVp4Ig/zGTE3qY6p3Xc
wRhWe9HKydEONQ30Di2zURdMZw5vEcOSCBlsDegqMK6SW3oNN7NNzNC+UkAAMjkK
Vnbg43Mpgt06c36+9vzmNwyO/6v8RmbH9Oe08K14UW53FrUb+qZT35xSXYYD7w2M
7ZgqgM5/vNcHT+0jAq8mWHDRCjEaa2J67iq+BroyC4t8xW989hicjUvJyi1rros+
TA4sSxjFh3+71Xt7o9Lj7HaDSP826xoBzks8ULFYn3fjom2Gsay2X9XTNvoX7rTt
F8u7SROb69OuraAQpUNrV1ykfGvNPZ/DJ9r/BE2UPyQdspHW8m7EWFxIoR9/bfgX
SZX5HBmrwVcmxKkIztUgka8v32/O6exVfSH8qWbbeGgwd3qXgZAMO9ITx00cLI39
WUfGPt4X9Pyc9bgN+qZVeSOq5GLd7VsfW61HT8ZRdqjLd6U4Q6EprNNcQLx0GafG
B7Y3oNZueCblVlG/QfsfKNwx3eTikNyIwO6AXs/Licf4KDze7gFYfvxL+IdtwTie
Eg6R3XtId9Um7ZG0PTFPvLYYyIpHVzBY6wABEMtcnOu3H+/H3zAI1FFfeREswwi/
Yho5/rZf7s7f5DR85Z9H9sRjy3s0Y7pGADWpruWDSmsgqIGaVJFEmrEnV+lw9baT
TaZyEC/0OQoY5Pf7gstl8/Zugr3f+oc7AUYbxUrPwQHkmPITKh/jN1+ETWPjdsaF
NxYXcy4fLQMLqb3dGMtZ4lKhSBRsWYgzlmtw19MaHdaiRZOR5mkBYQqRuDQ2mJwO
O9PiUM+6HcmC1PZUHvU5HeqiDHCmd6sbcI59c2VCIjJsdvKswSMmQE0rmAGpuCtc
e+76AHRuQV56ZMaFBkAdrPWSXBLPinfsnka0wvUQFDI/jI8Zbe7DEXW33rgRcsBg
vOw9g5GMrWiAGnfH2bzIIaKFudjA/3EsJ10rCD6RwERAlIQdK8nQUAA0hVa0UYqc
4NdCtOnl8kIXDf8L5e5wHX1dLbEMZ+oORxtovki3gP3et6C1IHHwXmYtOyDu/J2e
OiSbphAHYC0M7PVGNS1fMHlzRFuldjwDZbyRMhZr1VDsaGS9aegw2B+gfYFdZX3Q
VGtdvyp2I+jJ73Ts5Wx1dISWDKkjnj//aHnL+k0BYr3VCBqmm4AMkiQZQfCk4+yh
5ie6TsR8Axp6SPToQkHW3BT2tuybmxT2VYpt4M5stYlNI9waU92xh5X/c91dFYHA
hf4AWA5WT5k1lnSPVC9ELdNb03qRue5Cfbjb9ETBlO0u+xuz2F38IrH1C/XUMo/J
GYPSNMABASuvu6ejpOljSP54yzaCwKoO6H6Refj/tkmSCJn95vCwL94nMret+LjM
t17VDYgI3wtD6k0PBwcLFp8E6dCHld4SkJV5mD3diAX9pNZncxyON2/PaSrXEvMZ
3E1bYEHXclqeal369gwGYmU8qem/tTjdnmoRm/le1vhnyppgIWvs/taz86WF/kwy
YZxixMHAdsDU332tN2wT3UOVAvAOk8vRhJrcIAj6D4xadbLBdMqShWpjBBandYwD
rcgzAnUXr/WnuHlfZVOjvig0km008wLBq9juo+vGU/D6wwKy3sUw0rQyNMAyGd9S
g/n5JWHnG4X1yO6s01BBSvi78I4TnuZIjV3IMdX5BYdSmXTeepTwJj1f9qFyDwX8
bGMN7jL1bjqW2UdKVZwFI6eDLTBnCCDcCRmZy4Q2X0sTqL4mogurx8M4kGldyeAn
b+8kOEvYQpBnxBq5+NGVV8OMmFW+SvqTzHqHaHfwfSfkVOjrk8S66KFHmEz0gHEP
2FbTVL8q0i/5YhOwZ+eye7uYdqCjFdP2xqiqcpVII+dXbDlpt+FtX1INGWLQvq8M
gjlvZHK8Tun4jBazOXWpjpbWr3yr6d5xHbZNhQGT44Cz6a5khYgpR37ns8i77tYB
VpcQXCnbZvvE4UyJwSVP69HZ+Vm6h83lTMyBCS1ayk1QFZlR0eaKY5iBtLVt3OpB
bqalQxS3ZugxV3BqTm94vcdkgh9/iZWznNj97vL/0pwplpAS4I09Pdx+rwkbKIoF
ZG1fR0g9KhEFjhWdu5tvkCpyPJkupqfNtbudQXjKapYpFl7J3r8X5QJi2JDTYO0N
6cCUkWznHM4/htlJayHTn4h/KeyixgNnYgvXrBq5dQyiDsDInO+048L5kCpv9aR3
6DcOn5tgIVgi7nf1g1TdTp+nXH/ypkUos2HJEWq7UUVAWUBcnowzDw/tFzwsuAeg
ivYJ7tnKFHojSlfXRFs9z9CSVe5rJ8Cp18cpUH2rsVV37EMaa9Y6PFj5I++nmSqt
/tYbg7PkUZ3paUtacaq6Y88AC6KUO2tODHcoAxKiGhF43w0NtCU4xhC3Pwo+pCBE
/lEQ8otYs5m/rih2Mwog2kgYUluEw1ka8Gn6dYYJ+sbeanExF+t9l6O+10Mg5KvQ
YJpFOXPRPNR4pRLLlInKdcgjEVVUYAzupO3KPUekFGGhfe79jMLeb2gt7xTjkSQk
gehYbZflNdkio9Y0UAS7fjBC/lJoOkGXOnwmdAqxQEgt5zAHX1lpCNKwSQifce05
sdFrv0bd5H1go7oDrVkUbr81P23rOobYYoMFhQmdyRW+QjjEU8xIKOeWqM468sSx
dEy4yWFsZWfeiWnMRmrJMUPhBE9WhX4u8sJCyeho0aAhHobIT9synuATLd1Nosx2
90TJqRuj1x1e6PG5/y8mDauK1hbg10qvT17PoTzIZvv1YRcd3/ZX2K7RVLz/5JaU
Y/pDAN6keE4Dd8pOA1Uj11X42LhwNeokiOeWb6RPVqRlUEpKzUbcHfC7g0e816c7
idHuzDV1D8s3YX1NyQuO2h36BIUZmtvUl5FsKtLbQg2r1/5YI0O3EZNvUT3rKff+
e4uJnSjKuInPygEbcV8wkxRRaYggB62cyZEprQj7uGy5idp6z6L1l16Kfh1M6vKO
IQBhdRexytuEU2WzKSDTLGcO2kDD6zMEmyPKgCAmJeT4oInUBd2Ewo/aOtC4aWiS
rXemCkgY5PV1z5ZIVY+0pR/u12IJH7UJC2yTmBofY4J4H2VhF9wvqUbdkRLsCum1
aw0s/b7jWv8+inlngNw7kOkn80f4AL49cOuWaUyhX+JkHJdXMSS1b1/FFkBXvHGL
mU642kO89gf3UIzRG3iqiLPc9+vWKvmUDPW41j/J/b/AmILxgD14ZQdQtuGIfyLf
PKXeBzrfooEBz26rTCVqsJWXDbaen8KQi5GYfL2tzX8BHQGtCpB/L1pqmUgQ/cCI
muFXqGw62t9M2DKjw5N9r+MmuN3kGz0a6W2HQ4KEAOoiHkayWchF4h6WboTl7U6Q
lVhjBYh5dFxPZ8xU/LlmbOkRVPNJMstGQ4i56TzTJNNHSzXOmQTcNjpRBYnkcM64
L9qhbLddYkhRwKmGgKYO5W4jsFD0mgjRZNNd0+AuCZxncgO624sNacx/C/01kEEf
KcdMzp1hiyngZSakUpZ51RJfWXDTUR93SDmmuL932KVYhywdLxm9tkmWbxYKvw+Z
F+Td15vWWFTs7HpBfq/n6scbgvAzPkTc8j7quNWw8aQqSvZ3u0grSiHZ7N2yAPAc
IGihP9Nlz8+a1oqMouYPY1EDLCPKegDcA47i8Oyb3v2ehdy2ydfE8HQrqWIPASX4
4W300UHK5/CAJl3Rg6qsvHCyIopzqmJWLLh2B5J717Sn5TicAegar2GpL3C8J39W
SAfQPwfQuvSUNYRaJ5+u32NQ/M5XHduW1tICTIqIiMD9KZVo+UPiZMC4fMLfI3vi
EN0x0i4s/x0beYlkL62WmGsLpV5WbafkX0qyxjGNlVy9VYG3cdslRmKhWyECEJlQ
BPJq+RfrLvWv1i/sqyDELmXy+rCAcmuQkQv9rMnXAVWKHkXlAzEkwxsPNietKw+Q
m/vqm1EGfOlSWuclDmi5koeCpQRgc8k6yodE/NFXEcGRdzMhzGX6+w18xYj6siUO
IKegnJ5XBuzTWGVX33tCFJrNL3FVdXzyriW4dU/+LrcvBqI1JhIr0dl7mqaqdLCx
63a/QjjxFi4KZozUIggrL/GTQE4ntNaq6SnOteEJPVn39snsXViLJWjRpUZ+FGxq
Dtqo4Z/w/6nOy04B60CzCrDUC3mgMY4/OGifq6OL1k3BKgJTlB98ecLLwHYxXWw+
k109ZOH72yuuGG1lErUs+ngA4cTyENBqDAV/Dh/+NLgJsP7Uy49MK0dvL6xaeacM
is1mz6Kz3+EZYzFTDnfvce8edrfZ3Mvkc4YjC87zhIkkwvDv0+77Npdi0EMxAu1S
FeiUgHDrtlQ111Ml7JdKA+x/DnKlYStP4Uc/b7uQGHkNwCehy7U5JsFBZdOnddJw
o6689ff4lLxp47z4fDG1vvFwv5r7iqkBp+2RbitQ1Kh5xjlSZ5Js55RpZ09nEIGI
8hVvKc4JL8F0U5YVnbDb2nAqssnXu3pAE4byK6tZn1ipvuXey0RDA4Op0Ji29gkt
SknqZ78RxWq/GQNw+6lSwFLoW6FGCQshG55Z1lthw03WShR+U7rtonVnOZB1N2mi
Ooce1u9g6NbNgt94Knhd73ci+G4VRF6w+HSk+jCdPqsS+pBCOny2wDFoBPqt+5kJ
bXkXsSLj14uDNEHAs8st3TZ3wfCJKWMIfWzLfqXV78J5DTRlAUufp4HO01tK3Flt
ugkZfHnjGWCSGyVP6gmFCbaIln8NL7ITEvy8vmEUoq5OyH9ArpMrcwhHDY0QK0du
EbxyGoSgxM4FXP9l7KEWItkJYhFrR3Zi7gmrIqL7rvEEy52NJlSwMBsCxOjNqaV9
D740HRdyeNObvkm5SdZ7meHxCf61/nAcVt9K0zSni2mSZPO3eXOAlMmN/tnkv+Fm
oWtxoO6HV1S+3R6Zdt3an9Cs8aq7YeiYMo5IbgQo3EXCg+VYIfEf5ZXvc9M/CVpN
f6/T5ZAyAQsuN6PYAc0ywprCgB8lv0L9RAfIbTz3TUNZ1avWKZO8lWHcnAWv+GXr
vAS5Ulc6cmdMcp5u+z+5qougJs05F7Dvl11mzGacVVLZVlKjCDMzb+psWWsPB7TI
zow+J7ICUP+42kKLNn9+8V84LviX+fpkJ+C81SD6CZjxWCKK4RpVGW99saZ/Mw7O
nlo/zfdQe8Iv5OhBJlO3DqIfhttfW8yDhYegAMvMhwJCliPbkEnFELh40JhHjqtu
HE1HIxd8ojcuyn7MPgAta4dDDt1sBbax1C4CiUhjAkJrRMEKEcEthoUNTEXaIeIG
g2NbdQ8cHsyJKz0QuKAiFzZFVJNQGnRw5ckXAwS+0LD9EqwjKzW9ZqTqz1SsymA0
h+FgNX/VvuNeRgv/1abiKUDmT4umP431ETsBRCVlXdW1h18gXRjpviLJRUkNhOhE
G5ZRmvh98xUESXe11Da8SF/jEk8FJUJPyzxZvmy7oINNAZQm/dsUF1UXZUl3Kx+p
AWnIWlPRlNvWoIZOK2zWdkSoRdee9gSZ7jhQTV6PZL0tM5ikASP7szC6+pQqa3PX
xcUby8ynLqGNrSbqrjcw7qFWvQYHsm85kw3PkqahC6rll6PtXnvdMMzt941KrCZJ
CfVB/QyRDSNZ46lXlbYvcajPj3w2f9sbKADnCs/pB3I8SGtCqzD0IfTd0Oayz/SH
bHnQSSdjShkRm/Etd7RNxknD0/RJRJnZqO8R3Hn6WsLJNSSyOg63A87/+D++BMLr
NnwWNZpdonkWExlMIAQIVXc/dj/BwotVhDbyrxMlf5ysVlfqRqXO5W/t984h9VpG
syum5ku3LS9Kcbkk5tk9+CmeAKDCUOkNXhF2O09nOpDcW4Itu8e5e9kJ/p+CgCVt
2gmoFA7sdL7BRUNDhc3Q7CLBBc56FKftRv5JvzmiLdF5YJTrJYbJKdVyYtWdl7sL
nBP/YIiU/VB6TLEUvTSxVBaMFEy9AhpO0+x1LIOY0oSzizXLx++y4OYLxr2Upuxv
1YatGCZGXgkZDrZA+mJow2iqrpfZPn+YojQZlI0blBfnGp+jZc4weLh+DoMTd5WX
6cvW5D4dbJrEunZhyUB9gDSP71apHuscmXkxwjXR/lq30CfiewFpO9jMNW1xzK7R
0XMGg7GonxC2qCmeUZ0yAJsYOfDx1sxUkq1dniYGE9pYYsnrO5sRG4EFxDMOFBSD
cjKqg/9KH0BcgyfUpiM3eLon0lrIW3IQQGgChoEAjtlc6HHDAX3F4yp8xl/txQA5
TRXzHFJ3zBIO79ANi8oloLap0F3zuqFeqCmJ4C1BIjPgKy8ect8LXMeTGPdy/d7v
q67LjmZZb/TFMkFmmOqiMfZWYSFGnU68tGaamnhPYvKb0oDJL0DNR3Vqk1z4CP4k
4SXepVKLoC00Q6CERbs9L3iOKatQtqD9mEcB1qz+b7IMYCZa+CQovDr6rULMrBO3
Bn4Q8iyFBhlCgkCnK9QvTsqKFwkV21W0UsZVmxQ2xXpKmp5KLIyiTKakw7KDQlEe
jDUXMkJBMtIPpNmKcEdBRpyme80MYkR38lDKqtNA1egbgpxiflM7QnglgDCHX5x9
SKHG9Oc8ZL6FbPGsh0KJTcVbPZgc+WW86YrLx5SEoXeiGEeRalkXFc37eiL3hzyc
gTRyXcxMAU3emHfpQTjjWU7SYbjNSwil4nNnnaspVbhc39oMb3HQwCKTqgIMCVHi
c3ZJ9E7uR4ZME6sSFKpkYw4mviCH0YLDLnZ12m/T2mU2PmrpaUrdNquKdZ+dHKmQ
FMi4Oe3ZJu4G+tY+w2cZwUgafEMTM5VjNL/APrmXvwCv99ADH5Ym2rJWOIlj+cOg
U2qvfTq5+i7oEp40kbDcTZojU90XOqCXzaAXkCAwn2orqxuXllkuioT8Mb/eMwFK
VasBIIY3/+LB1xOVpIFZWcuGE81QQ2h2ugdqnIIk0Lb9LTLwSmb+NMIRRo/cv4By
Q0aXIVsSej+El2Xq8kgvcj9FqUgPD3EsY/gEvBI9qrZGp1oDAT3Zg69ycEA2ezrg
VMyOpU0bITcWnqPklP+boUw0ojzbcDg9l2X1V+iEmzr4GW9lJQ5gNGbQkfHouxhQ
42+3qhuSZbq+ycXYA6njFytFCGvD/UTwP/KYB90Vc0296Cqdrz5jNr9bJJOZLQVF
j4RfafGMcsPRog6iKsuDfPwPCP3rNpGiAqU56qFARdxl8qoYxODaaSswb8hpENTO
uuTyFRJO/B2ANICfBWKFvJtEVWLO+PtSYt1HoXX4t7cvYMdQoIrpl7VJ7PFht1b8
vTWlluRQtWuu3m2T2AorpcnJxDUksjhp57Y1ncgFobCfL1lS9VmzU0E06tD6ydzT
8X3esk86OX2qRQ4hW90UzGfjgs9Iwohp3ilr4ytGi+y0MtdOlAlY/Eez7ra9oaPP
arQR5QeaFsv9gVeZDsheag7I5bKRJ+2jr7iMRFYbh/JyqhfwsSPMz6YDvGfS2kHe
y7vZdjbQak/lLtSCs2PU9VqW8IMUriuWu21vyGZduSmtBhLQ+ZOmW5zol7D54e6g
iOocRdKV5nZV+HQ1TqD2TWz9fn3jWSlqV2Pcz0jazW3oVMq/vovUwSJffG7JTOnV
ZEa+MRN428+NaFkhqrBHK/0zjPSJ02CPxhCCWVJ9ZHXpxxo8z6JrHV1dWYlNXGS+
59MlyxrpdgJ8CqWxu6OYlepz9pjKPw1Wg+LJ1jOEDVikl2XPaNz6zUKutpbZtDwV
E7i9SUBhMkBqoeX7Dmyxy9GKyJvyIpZNmdVtDqwvlr6DrDjRID7tpZIhfs/6H8Ov
9KLlnK1SBtwvmxX3cSN39X5eRD1+FF3sItFlGFfTKGe5dg5rz5JJB9+ElXkHWrtI
YJR0muvdKqVtvUeALV9l0CT1PK1ovbk0iqq0RnBBM0RF98uphJ85m+HBLahE6Tlc
Q1tOp7tyQPdeRLGFM0SPSTf0Tv0rh2sNJuje8aLHRwhZjd7xVoRia7/xqfS0DAw3
eYlYMxMQTedvsOWS6ajXCEKVzd3ZTJVBzv7FTJcptGe8mZSqDbZsV4HvoibavaRg
QPlas4EYvmNbEC0lwtMOOV1vUfRSMYrweoFDtXaaDWzVrAaxUMU3ChSGVGGlvCoq
rmbx0EKbs9b3DwCBYWiNQPoe4Ao5Jb74PsQ2+njXkdsq4oa0oUQqPKxctNWquZfY
kzXZLWSSLLSS1Q38symmM5wcmiR1dh0iFi8v+rpkJE8xlWipFU5wEFftn63ffKfk
0Un4WhnUdieK+bJS4UZBCFAbGDaiDj64HHXX/mHPzBNgY2nltx4TLy3CChG8ZqVT
D+1vUcwoLD+Ir2r0JI39al8zb8y8JOV3SgbpYBltBU9r4ohO+tLuMR17IXSZ3rT5
yWZe7b7Z0SeDceizcdb/rjOxfyyL6/mRJ3dWzjRJHN9rmv20pT85yuws0zoVC7cR
GsDsgtAwzpXTYY7L1oA5hXW0t7DRhsT/OUi5sC2wahM34AYMrFeaE/DWAGetLmt2
HMu67UfwvOIQsLqHOXVQCgyS4MHHrvj8NwMUK8vcTMCkXORDuoPxhXR8xvxq2HSh
LPsYTZpdTu0CUdtXEZpfcFZuvanEDXH1+bMPbhDzONXav21DAFurKGoPr87ujbWK
tB2slC8i3Bvc6KMigmNjb3qYB/5a+YG3JhUuvEFtbqdIPsSRW1xmmTxGGONyl8Jn
9rVMvBXkir0CLut79ms/Eiwkomk00XMXA33XsjPLvE4IlEm10SmkE/p6K5tzxiEq
54zSbnwZrFPGRPFJhL5q5w9MVYByov3FlZARyAlAxCniiKAc3ivE6kNUkMW3n+bc
R5A4caEgAi5zMkvowfHmUnouQiZtULV1eEon/aZFfA4d9nBM0STLQevmx46IckO6
8ZUXPVO0+4cR0tnuDimVIYAjcDYtc3AklojxYJbqMPdLpB0jQeZUtDCYdHUujSbH
JHJ8ScCF8nxBkMNu0BqYhJOyD75FtL1yqi0VGRFthyJrCe+avwKdAkpgHVfmMnnv
5K3mf7cpLa5F0fpgVafDk1bNdVf9aL2rfL1cgPiMIRGXOvnV5/hg71SyLkprZpZP
S75lGpn2eyK5cn2wd3OmcUwxVLyxuH8sDGDk2YyxWu6uMK8/bke7ZGV2jApQQ96Q
GgmjFjEVGwGznQvTFSvitczR0dlrNzgnhlqj39dQVY1ioizo2Q5XSO3Obl7Chzro
vmng7Amlx0UAdX9oCyji3RBt4lrrkumf3sEMs52BeVzSmDs4yqREdchMNM3waIyR
u7f7wlo8heY14efJBdO3zMSauBasYFzU6iWViHeDF6tKxqMqArDrkp9KHq8xQAfr
/YO1tu9Xt7ga0eWM5vATMHXkxbXm02WFUeYd6TPfWMm+nxElACHVeNpF33JbjGQu
ufT/nIAOzbk0swz0Sok1PsSqxNjgej+3MQBqp+hleBeIvQ0TwsLUtvrPFlncLnSe
I/qpHp7Z6flWvkBKxkIsRuVh2jmjW4/lbgtTFdsiHBezXCJCkQoe+mdIwbYlmNFM
8qAEGX2ZraBeoJnSPWb5Lb16jjhTCYt770obcRbcQ8oGfXD0SagzpnS3sMyRF9Ab
BfRUPYuMCoRrl0IAjmYiQb3tE5Uy2oUq8kTbkII6t2w7Nu0D4gkc4yWMCkX9GN+H
WXzkXyaJJePLPn7Du4rLAILy3Hh6+0TJzRLUIHFD98wnwxcRRPQXpB0u3gd1K1MC
O304CAoQIzxO14PM6KyJi47KW0NYNirqLbiOTFB+M2L3NPYxsAk53aML5SxkoB6C
Uzzp/1WK8HtLr09ARqYT3WqEp0p51i6zaFXcxPUuXR6WRkjtakxT0joLArVEx34Z
nRhk7BubgF1Pb2lkKNQXyVJNnUcuka7QdPEvCjgkxSjuaWUsnCmcwC1/wq7aCmDr
6+wv7LiopLUjFryHxw9r6I5/s7Os7bf0wAl84e1vdm/0SiHoLAJSBz1RRV+VsRaJ
O3OL8hBAmjPhTFkCinUyEDQYzTkJ3NKcr+E3ZzbLOjld2UFbE8Jrlt1t12aGnunC
kOMdsPeBLDmUKHHZXK3ROhU1vuGXYx3SGV/P/QIfQfCPpE4Imos0hZ7V7Ryl/iG2
v8hM/UG9CbYaBdrXMPKo9eEmynPJZ7X1c4zDzGf+YoPLlvXMJqOqW61L+xozL+FL
w6X7d4ogm03j4QSAQYyynIP0PV6l9L0XUlTT4mrUcp9z76AQP3UoWZRxnOopOW0J
g/6zpKYre6fRpmW0cFCbrtMZM1mM00zdzcwr3S49p6xEKZjYYlXnUIcpZtOR/UL8
oSL8QR7irFttmWWxguCzAc9syE9ZQUtuUz2n2CUzEdpJLRV0lGg/PssC6JTCU/kd
rN/jOwQ0kwJwn+ptVtrgYdyk9fxY4PpkAovYqxzej+Dd5ODxqW1ZVVxaIbHAEene
yorB5V2Ogymb+/yf4/5vBpM/mpe10cJWfvys13UdGkwH2xkI7Btq4anU0bP4NNO/
PWLZ9Ikf6n8V6R+GSVTaBG9nUd7F+23SBYyN75jMrV41grGkYSD7NnqXpaMDPkUT
q3uYmkMZzvsBCf8rOC5KP1XsuRynrDN5x252SX9v7o5NXiOm2Cc2m+RZDP/Ew5U9
E7ri/ulL4rr+RYg5nK6N6b/hyeJyvQrkQivwhJjioeHY+JsANcyjHGDKAq3DLF1p
myNYvLRP0hrhd0CbRJw8gGPb5gplNuTIcodArHJOmg5w60p7inhROi0NaPOvV8Hu
3DM8aXRs29aof3J69SOtjEvUIH4Op0ewNTRnbyWCK3YF7HDd30JDqnr9Nf3d8yNH
PLcFeZAyN3RDPuoqscuv0YZD4mcwYyVGrChApNNklSqAENHn+5/tATLlh0z7BJL7
eGQbJXpCVC0BuuIz3W+0NHtExP9nUu5mICcDAQ0rvmtSVEibcW/jLCZZ2U44RSZE
N04GQrsl92lFvHnZI2V5e2AeYYj4sv7yE2diyy90X86jq2756kCCwj2N6tIrOwMK
2R+3XGLw/cpDpO1kOqfzBU6fMqnDVEL4tYuBVCELnRHgCEGmQZ3AhVSC4NPNRBKW
RZGthjan2u8RjVxvKEPLLw3ZjgYi7VsvzxUrid44FqfjO0Uog2J0Nw/XHkyMKBGz
6ITxXoKJnUEH4z4//SU1PzpkCvkZOsdprBDw/9wSLa5yK648J7pPyTckmVE0E+B9
rHSsghvO9b88k8F01hzgm1ugAmeChOQBa6fR+f6xksQPgR1OCWFRvmKcCmPYmhcW
CKCDYRWCaYa/j8OLEsHGN9eGjyc+LBwYmPkwSk1lcs4i9X0w9BCwmk955RXoiTfQ
3zO4eTHmTheO71XUAqKU4Fbhv7lW+2G7zfQfil3QBVw1sNKEIpYoCh1ufTHabu6b
444pJakDU/7I4Di7Fq+GxjabRuNajc3N2O+7SclIirJmTjXghmlkpvo6dXB2RNGL
JzsTLz/ErgL3D4rTKkGqy78oHA50VFUCos+ZThM9kUX4SVK9o9c5GeM0Hjt5EXxd
oxn3c/1LKVaqpWhFuLtD33iGvFgGjV1zIafXoU3DPmhstU/Ke7Spvta/LGxAsAbr
0nGCWxpMM5tytmZcQFfQWBtGs0WknuJlDhvbmyEPuctiCOJVm8EuDT/aB/SQZbdN
kVWDx9YIqaychc5O4iCUQliE/OJscKAkQml1QyH1JXFdaBh9HZn52Quc80UZYLoU
iiOJrBZS9e/SdSwe+rY7ypD5Y6bLniLR3697shJWMPkVo1y5fAWvTzeCwHJrJJpl
9fffq9ITJ0MhiCvD0XuqNdZVVqtLXD4fXgwhS8j9i7Lvxabe/uXnTNpgVjZ9PiPm
tY25Srv9NgyZKDu4SxCWz/+9fd25RSQzL6zrheiuATnFBaTVOr0Nt+d9XKnNdjbR
ehu0v12oBvWtgWoNH6ngJzQceMXVXWYBuXjpjIDpyqKNhUfu2s363eDp4hCxsWcC
ynZYWRwxImF2H4kVZKaVGJ0F+RTiI1exRAVdOBzMdkF1y3QOjGLhUCxaXeo9lse0
vH3wIWxIrXXK2jiCtoJVAEEj0n8JO326tp0CDabNsq+4vJZ7v75qql84m04JAiVh
ihUN/NYZ5ao5jIqhXrXbZVIXetpyzMBFS40nhi8CbJL4Bzz9ydfnFJpDiIB6Tilw
UXyzLedt2ykLl8WM5zesdepj1hU/uoqH622UqikBrdEBQsgQVgUiUy1hRBb/15LE
xJH5zjUW9//qS2Xb5460T1K0i/RkthCgUPjTVYc8f42DtqDtlvXTPEeQ8qJfKhSF
y5nassiClGuhkJMsNJbQAACrw6YAyE1torMaFX7SBIJH/TJMMVC3j4iO5Bj3TCAR
R2I6EZkE2Y+K7wow0u1p1yQCh5MYuWftFUDTkED01RIgmMLCW9iHdzfPviZ1ZDFP
0++OJ55x8YvC2Uj+Tpz3cs2qWgPHOsfbGqwT5z2sb4hzWrUA4TPTe5l28NjLM1d7
ntlzxs3EE/BJQy1RqRpyS9AritaM01Y6rscNdR7KTNa8zAzZ2ufznkkg/gn1lAJq
Ge1o5HSHILrs1TOe/towYB+cLEOzRLQ0XhkTeWK14S72hX9HEgJI9fmm5QbzwmC5
UYmVqBHBrJDhAN9D50qvQ7pB/bMi3heTqYRi4GV604qRKRmieLbFj2i/x4VWQWfh
QugTB/Y79Oqot3HzJcMYxf/uLm8H4ScmDSXI+qmENhzm9DO44c9YpzPadeiukgUt
9bVUhQnRLy2ITerfm965nrEhOVWmc22OtttRICZAXv96QojPmXatr8nkF2K75NvJ
n0W5OrStBRjWwesGhs+3pbsb9eWG7D1OZlb8Rqh6SjNrFgivHxnKWFpTrL0+P4Es
6TIZihmFoS99EpxeVOYVJt2Sn2CXJ1xahXSkkthHPUUpIJkqR46AeNoQbb+FtLDp
jYnvKEjQsZEpYGNHpFa/XufTPbOKsi1sDqZhQDTzdFQWWy4vBuXEOs0mp4u6u6vC
N6HL4TMs6WDZF8oYiFBllJzBT0mBIraw8e785lglqjzv/+f51fkG31ZtZ0YO7OLi
KCZviTkui2bKrl4pIV1aFTLa5fsLAx79bK6u6kjXGExWnFk+xGQuNq7Klg59pH4Y
AeYUWmOELGrW80PhJhYNV/96gZEAioIPjM8GsIxsHLiXXI8Dj1VbmlDLGRRqneHG
zZHh12sYDsuoSvNw0xjBn6hX7Kzm5jGtH0bYrgNUyoRx54SEdqbl/VJ3CbJ5L1r5
xIFHTRjh4M2ZVkoL0ucC2Tz4g+BCuz7BqzBfPe7MclOs8nhl8cV8uMyvBdSdrvG+
Y2l8JlZ898hrW2OjFrFRValBCUa6Eh8ZqKmh9EhSa17FXVKFk0fvu2Zh8gMXtG4l
dJNGfxmKSbKp4/Cu51J47xhJ/1a5uiHB4vpOe6P6ik8+tokkcJQUp24fmhGHHvpa
bdrOFnTrpfRBI69n9Icgju8kLmkU9vfDn4gDg6Xa2Qsv+1uOgt+M2COzdkdA04G9
ecUtypY1YfeSyY5//d8uaq/SDWHeBAZxB8S86/1yn8S/xWjwVD68Rx8zuZuomqQp
bl8Ff3JlCvU1+ANNwdtTgODLzZrvzm/Et8AYlZSNesDhGvnsjnIHXuNF6BgEuIOc
y0h1Hl6APxyj5GSJ0v/PlYUEZIfrGG1E5mwyui2FSJYWTwgu1eMlksTYVfESssyO
tXXSuPTxCnrUfziSsS2Xp9l8SVhqn9p1xHwbwyZpiimgCQ94oaFNNcYQjmrdrICd
zTOz8O6g42BbKmUf+6QNk4r7cGXQxt5wvFtysOvQC/whcr7/8XxvqpErCIbzhn6A
Xe76NEKIBQB/lCubCLffBADICZ+7fQzCZp8E3CW4KDCPfXdkBZIGsbYxGt/ZRp5Y
jFPORl49P2yMv9f3+m7frUsD/olq3N12WfI2s7FGAdgRJH19u+SHwoGPCdET9lk6
GovbzCeaJFlTY0hSRoSGTMH+rQiiGp8SLRPkxU4WZv6N6qvvRirlZvP/a+908pHg
3FjRoQcBKsam3j3hofKZh0/I/Eht3bUkbVWVtKVZa2Hc3FoE6smf+eLYprFbqltd
ILoGIhSSteUmtgIgeRLW8YUlosPv+154xeU7EXZl1llzI4qPKH/3UfhEtZObeakS
r+arziDfZ7adeDwfRqbEWr7FrDABpOjF82Iqd9oOvIuK5uAFXxcvY8eaaba84/Ki
v0ELMNdfyvzNray3dEI3g5Z3Z/fcdPVeoAzSYaGFaR9mk5yOX8l1IrWZbc5anmbt
dHX6L7ROtnfxsoB85eNN+wtLsZjA1shuKAmRa2ZyYiDxNMPclFyppUgJdLrYPYhA
EGC2Bd+3E3xkro+6KvqVybT827xvRODex4xrQiQbs7OQ10T37wPBy8EGVGxMSE1f
g/DJHHxYaagPq7FrXzD2bSF6FnURDl7wOGNAcEQSWrOnLbp5wU4aGQDKv6B+8rY0
L69OOj6DAPMH+05w33DNhfPNXzF4MIG3I0pJ5+U7TWAZihuQTSRTuuhG+U1E/D7m
HH3a7XY25A6Jmt4JC65UIb9Tz5zYheahhCSYK3BOM962A1qDIfpYTAPZrupQZXJO
6o+SUDTxVLs+0jc8CAWmhi7dyyibc3SqstAZ6gVApm8BwEsV+BkHRteZr7n9IavV
G/Nirxjkf5wjo0pJOqWmOTge/7czsrxQXj1wD6KP/A/xxLIXjwbr9Nf7rCk/tucF
x1DG8zl5/mTqwadpU7KpvCfuC1x1B+j7lKSg0LwUJCuo4Mf09mJLs/8BqEUBKNDu
JMtkf+jjZCG/cHHqquXTozSa+bgrXMEMrOm/nkPGhpsKvPf8dIMa/npeI83m8s/i
vier651ljB/V44I9f/31hpdXGgXlgbMPvfXfKVKMdWcFAGKbLKU9DihrMBy5+fU4
SFJsDG8qiRz/X4bwP+MUrBAcBJt9FYVKSzwsPrMQ39nBIIA6Wry68MT4zTCkp4lD
4EF9JOj16qujLzP597Dk8CNZPjYm+vt1uOVgUiqXX0YksB5BcNwiWlD8FEuJ+yLF
HC6qChJI4qRTU7o8L4Gv90vKHZQCu/m4AXkGQftCp20OkhDGtErKp82NkseUAN99
U3/i4Yn5kqLflpLn48xsifGwDU5Np2hJFWM3EcLK6XTXsvp5ip2ji61uoprFLiav
u/OIOZCc2f+kDJgca46A/G4MUpr7JIgmPVE/TAGvvXCwzKo2Yrdskv07wkp0xqq1
wDYNYxl2VJlWCZHBOVM6t4SJ6CyDbdljEsR44PRA0EkFV7ZjkVBZSCb90PVjxP19
g0uxiA5prRMpenveBr1OoPq2VZ3yg9By36bgBiy8/n0OwxL0kGr3o6WTXsqj+nGI
Lf/zUN+8gkcKi8K93oGRt33dN54QA/QrVQBCnkkFJIdFIRppX7DdP6LwkINzZi0N
bD5Yk91UgSM82g2OrXjt/GN7/r569oi6pJggXe2j+2V9GIYD6tN+MatQ94mNoxcp
ltAV/fZUbNfZ27sJ02R8hh45DMdqr8IrSWL2S+mG9G7cEX10SlocmtE4qE2JBmSS
KCmAAGh2DCWrH8XRSN0XAXq9DPNWvy9z+hgiOTkZD5OKJwjzlVZNdhHQdlQCmteP
YrIsc3gozizNzzWXLLVO++d8EPCAfVbYGipI8XdVemfRIYx9XYmls4ptiRwwXtdA
ToJR/OC3xn1p9UffsKZ5zOklKNcAYdLnaivc++Bybc4TtD+g/Vlgg9/yq8DAPh/9
4GRLcihxMisuiIeWqI4Gt6T0M2p74JUeMZi63voYdm/8mqMwwy6ZC+OfXeC4tHdC
CKxpfDl+Wxol5z8516S9A8kKGIi3F8b+5IQKPmGgkkvxzuZX/JvlPyj6kpFU6/MA
cGPPo7lWLvdLYXq4SfZPgbf2llYBtr18+XFXzFGHdk0VpB6ORqOYuGwnrMg8A4aV
tfb7WtWKpL1w5JfijB7EjWu/Vbn36rwKglAItelw+Kg25hxorXjR8OA7EDIkJw3j
5kF5PpDBbbtSI1yJEt2JLJWCYhjWr0shLCTzB8ahqi+Sw5bwbrSCKf2LjzCePSQs
+bsMCxBJ3BNGPfsz+eaA9BxrOJwZ9Rmu4YFBWShVTKzkXKqgEHR+jMEYUm6Wsj7G
jYpmZh5ftyIYtiRqrK+VhkixTNuA9cGXsR1I/tkI6IdRfmxV/SgDE57slORNAmfV
NQQE2gaCE0v/L6IuVa/JwwTKVbDSPYMD/0NX6ghpSYW5StfLDO+L8WmcAMcySUhW
W4dqVddxkGDyUbj/TNmZaYMuaLxUykYRSwE5tDgyoK6d+6nQXYo8z0W9bKeuDCYe
SUyVMBb0qFBHDMV4bIM7sjM5pvythw40vTNxSbyWDaufvhtWb40vPXGut0vgSE85
9kItdujTrRgzsyMKbff1rbCjx/UEM3l3WX0bVC3BuBdjIJpm31ZElSJYpL3u8+ku
Zaoh6/xpZWDpLQRVzwKgIfXbj2djqtmQGF4CULf38xigAho2pNl1fDS1+GN1vRjs
MOevQKViEzZ2OSmUsHkeYaQUZdtAk1nDvvxQuSKBXXF0XVd+DvmsDlas1ZDXBTxd
Fp3h1i5/O59kKmuJowejaMvJT7zH28S859KDBk86gt81sA8w8DcXuVj9A5LYZipB
D6ua5nAokeVg9l3/TJiKtGmlLbSmtmO5FzsgldeUS91jL2OmQcuMiXL5Vbw/pNZR
5m7Ioh0fDN2U+lZOZB9v5OxyrFh/H9x0Ljz96ZkIhGvF80gfqYEk3EQuMO/29RXD
uYvbHJ8VATp6dmOEro+r+ei07Dup3xJ5na5pxPnZIsCbtvTNExShAvEBGRFBdNrX
F9MAkRq7BBz8bVOumCahZLF6mcUa/ouJoTUFQT4vX/1iuTD5+QPSOSe+5/FtGZbW
eSwdghOXpJu4OF7lOGZbCthk1HvCVTSyCF8DxgXFqlbjecNskmShgZX3yNIhPfKl
IEUxPnZJE6dPzZz2xaTSJOvFtj83L2bMLNioIEqG1mEt++mjym+eeOnXt86N7Gp6
E7NjvK7WSUqjc4Z6QF0rdCNlX+t4L9YaWiTsk2CVsjakqURwf5oRxDryJBRmXhKj
lM3SOsCTJHrpFWkHxB046z1bmceLLbTsmlWaN2JEA7zGuHh+JHbGiZs0bvBSMLYT
V/8Oj64+vsP9a53xgCHnu09Jby9FnZYIr3Nn9Ua3NGoSSLjeDHSqnDBaWTNkCr87
bb+3B+MKYSfF1czUgVzxNBsIHcKRMISEbEGrNv+7coertWTVaj+ki+wl1plewW0N
q/hVU4cx/wcnYSlvoAefnN8AIGrMwe0wJZbQy4AhiiH0t946+XUAnemHxwWIM5ng
EJT6/JuONOYH2gDMvU2jRPls5d5FoRzHdc9YdeCokY2p+j+np9dtZy4ie+HMA+9J
CEm/4vvAPt9fyXlbmnpTMSluNMW2TowoDk4jiDccvPLSv40mvIxQ68vT3nQf92WQ
NKK0J6Y+0r7i+73sqiy9vDFO6BPlc1ysj7nqM8JvlSfVnrJzrUOyhrUs59tn3c5B
MdGol8gVDAGIQGgzqLGNmFdAjBDRYKbgsrp75aqp7Dew4vrEA8LF8UB6q5YE63eY
8oefTeotZuhgdkV0TRx9Q9MN7TzOxXG0d25jCHBf/C8PJcvRsibk3JKffMAwIaAA
wDHyr/W9W7ynMatbFgXEp5O2ZQThOFPpuZc7Oqw+KBp7YAkdUIIctEKC+yLiL9gM
9Mr9kY4GqiXTnJ0PMsxOVBsEc4EJ5qGXMLuQvridaw91sBe/VBoiDN1oKPH0Gok8
Z/l9TjmObsYf2OhmqBl2oAef08lzbVWcOOgtotN1cKkDjLGHn9VKeYXPrJgANm2i
6zbA8AtWDtaLSIp7Xb+44XwGrPJnPICS1rQLY04pt8JZbjjGMHGOsmWbbFV9mByf
ppf3ln5jvdw+ilWR3FLWMLuKUJ0moKBsjBGKIEJR8fqkS+Ihq8xGh2pTt9q6h4ty
E4eoUiJ1+QjOKJXHl1H7TOsrnCbeQ1om2dahflyb5OAKVJL5//OwuJCGTkXoLheY
tbS9eUs0m6dKvotOyiuH/6rZzbJSYLY8aMNOaPmLF4wSqLBRNVqfTr7evx4KMVK0
8bsvwyOw42GyV8hBBkRpHyeXbVQPeOJAMko5XWg6yxpl+YcDLyz59k96nh2cDzhn
vAABGXaFdzP6A4PsHpnke/tLQAYj/FIZf3Ga0H469kNFqfElSRhxIbayDDOvPtcW
1Z0svFpyleAcvZ9OkbIhAmSlXqsA57URUHICIgEZsOhAuVHISDzpkRFpSjcGpHhi
Lku2DKkgsbe8eVuRvitU2j6ERcYxV+edXRO4orvDNTd9b9eZ+qLon60p7Lq8rmEw
PkK+PKdKCI9R/gfna3RC98Qok6khL5eR89KtMzX0IoLSk90OTV7STolnidVPB4Vs
ut4wR/fCUZZWxghQwX0n13RNVBcy13dhQrG81Bm2oZ+FImc2qBmTuYolF4qkjxMg
Zv3Zg+kNKXQe20MX06v604Kw5pC4ICEC2ZkekvCNeRKHin8mjcejXfn0N7mrs32O
/95y/V301cisqNj7Byuwazh8KPsm7WtvLJEHWjONkbuVphM8wkp7Cmi/ulhk/rGH
oC/+UePxAd0XUb01F2lJvoYgLVMgaZFo0AX/aNtS1Ns42CfUJmWirTuCV1EYOdX2
w+GxSY1ARymVqMXFarcqguSZsnoVjIVuo0tcNsiMoF/7GVHHQ47DNhpP+Rh5yJSn
er+5f8pkC8Zr5I4mU+C09meSNg7/x4IVk450ellZ+fsTPah8DFZt2+HhSUGs+cGg
kuLxCktTPq/MyAuxohf28ytd7/lSWiuTE3od8YNIdjLXS6V+FhLOGqj151tWPETS
K0Y43o8z8A0Cn522fTX/fhzEy9bX1qNQGV/YtzBMIrnT9Se1zhuR2SJpzTfoob+9
qXUHmUmKVRwMOmLLJjnxOBB9bV/m3CAJaJbtVougRuxrQX+2qU04/UJSlobXIe/g
1ca6rqRZr3sH+SDRsac85k1ULu6bq8OIfWS64xipadZ+zJJoAp3mUT+KL9PAgp4U
jnbJZZwpFQYOBCFxAnnpD7lSmqZEuY5ktjLtndQJU1SqZaNwhJCIkivEclFPMnSj
fhS2qQMKcvSeGuKJCQLv7kTMg76S+B0fql+GaqAuSFTj3adj53oz8awWtgX2g/vW
7bTfopOsi1524AJbfzaYZtHXOEWUBSFdBODXlkQ5Wx3CCff72Ms3tY6HlSaPaysX
iTkvujZth1j5cDQBLmrZNf4nnkfzppANa5WqcT7Jyyw0A2Hs/Y3o9HSbCblqp1hS
wUf+u9OKPeYO3VbRV3P/palkYrJP6QHGItAjqQh/Cs9V9u8clOE01udQI8pWSbCC
k2fLqR+fbwoV/KMKzPli/BPBJvTAybpXUpHAhojXKDlGT9kXnNGwe999hjoL0H6P
a8Y5Y/NOb3o9GvWw87ab6HiW/i3KOhGpmLH2dKfRHPOcjIiiRV+ATqzm3kJyYxJC
MD6XRPuo7dcqFE7JYsiVL4cpf13cKv6baaxOM/kdlQBaW9v6SunGRSfqBn0782pf
PtMRomFU5EYjG9w9GfcJlj/QqPFsR9LGcDWigsRwd4UALClI6+9bpvOgnY71Ym4K
RC8ab4ICaqU1KwTo7LvTzvOdfJUkNaOxLV1MAtxDvoj+yXdDTJrToDxA/oeQDAF0
Sy0mrij1IA+kUyRZRKV6C+3gSDrWk/Oh2YOy+21sYIS4XNrtGgDTBGoqR1nO/tT4
dngPwrW4zG4TWr9r5mj2GmSxUmLSry+ZcYwBQL4QgnRvfsxBsrR3XYIgs08EmNwZ
+zVTY/NE2LD05BIyoZKbGKfhgwpCJ2C5GnRWY4jeVa4xQ306ohdgTSdvwdfqX6B6
j06cFZbw0XoxeuUMEKQPUoRkvNBntn+TZzvETL7KVgQYG28HfR/6vix2Vd53HgX/
Lc6GGwfKnlD31XWdyMfI0dv1BXlZxSDxbs4eFuByQpKU7Lg3q8YqIM5XjsOdNSYH
RHIthvS971XcYnJASk8qllYhnY6dxW66Ayfj0HlcgensYmsiXlJrrCcMxW26O5ZA
1uTD9fDq1kZVp+LUNr0y8PZnSBTpcDRJu9eBSoUwtLGOYSqDOnGyQ9MRcm7/1LM9
c67wK6DhLLvGYF1l43VZjthgV7EeLDRkPu4LdHM78uPCZjTJHImv500VrMIpwn1s
Ud4PyhV6f3aUHqLla3LjJBlYMaCZRBvBOA57rLL3yxePiFGmtrvu5glyht5L0woe
ZGDsUKE0XFci/GJTAHXgJdD82iQoIX+ucmp5Cmr5jAhciqE6oREUCTXD3uYhn/pv
WErMUfnTkX9R3ooQ1SPmMUBhEg0vcP3n8BEcVzx6dxWFCZuSYM78SGDMzxbOqiYE
Mob+iyRG80wII4Zoo8AYnLsYenqLGSKlp4kSMQE59o4hyNrX1D+DOhxVyslqoTUU
C1cFcRzCgzXj8oeCoMlHqoNaJjQs8LQKUXN6EW/iQvhc0XIYc0EDngtE2roCxFT9
psbgnRCurHeC8fysfqBWg1gGSbMV67DM/VpeCIYPh3Cbwrhnf/08Ars+e2LlUVzr
JsXF3hif1uf2Tsc0aPxVPfOgqC0Luk/qgN4SpoCwZB8TwUDO14A9MvExqLgIy+84
cW4RAoRbJ1w3oHOuf6TZ8/mnRL/WZdPJZEdioLaOPgvh2U26dW/q7zc6Ubt0XRL3
auGb0n2j+zRwvYcoATfdznrAOSvos3UGJDd6GMWwJEfu36iCpsyYVXxGTFswMJtU
j6grYlnsIbm/IveqWelbD0xlzvunKvfQ0yjkS0Uleodaqo36I6KmNoJGbMSXZY/b
5Ttr3zaQJkJZlkcsom4DfjZ2hN8VqAyG8GuLPtp5+UFGuPCcuvuCJcZESaqnn0nW
EBZ38ag5UILHRgAJ8cp/QRO8tAwMf3MQMK843EK71RlSN0pa6ZwWVAjBXFDAO2V1
A3X4BNw5LGXjTHvTlsZWK2LbkVPMxWaTj9o2nXfPgIywnCvPdbiH/q/AABh8kr2B
8CTI3xpe7nZNBaZ4ZwQ6FxivXPpdtjugI82QMa19N8SHsBulBbsZXXwVqbDSWbrm
fDXKdklls79c7szJn9hPT6xjnvDEYcPU4j/HU8j6G9Nis6XaAY8m8xfIFn+M3eIn
mkQWmPDdzIlyyKyJSizjR81jSxd3akdkjySyq8oUq72bKiIqlKKe9pa+T7w9AjTv
QFi+ojzVqMQnPdeBr90J8FQ2RtjycloFkCTeU7QQliyUky8aaZ9ju0nm/n9sWIx/
I9wisesUzvYT3qaJHwI+LFIgZohSCBAOqUX3M06fGjQg7gKCohZiigC0+E5Rbq6y
30SFwHkGVfX1Tbt8p4l+pGfW3NO5VEmwtx5Yw+Ijv4TqHrUN/np/WedZcNFc8lGu
9kncHp11fj1OXlgC839tT/VUC2/hbwzTef7H0CAWoU7b15s4fx7EHeV/74Htnx3a
k5NsXrhIU0vJPHBjWLv2KVK1duhebw4xNrcO7bPOmu1PB325wGaMa3DS0zO0oqm5
0KhsMqsmfYGxGlsNm9njVyzwN1I8p5TVknLu9yxQuHIKx+JsfbRtxyguScpaa1VZ
D30S0k7Soi+3JOWuLepe7s9NuLNqkMHFtPdCupccWAqDU0xaQQu5qExT2GvoCGQl
IN9lxsUccQw6V44uba9zE1ASTjLsD78rRMnIsoUCfNa3Yl2HWuUBecF+x3ckKpRM
lcRRKyi7l+NuS2Pioa/WAyjfuNhmYFCvpnNlPoIfncAtHdnwiOH1vxtcAwLVjHM3
2BRq6YLRDc6bL9mG33r4CEMztR4+ciKVDjNmjXH5BOWfb3G3SlEu+5RhFR2bJEeD
p+eDshRY1pfSJonOZR+oP6vBWnKlwlMRBBUsSbhEcn1WXExW9GS3JzxWuyRoypft
2GLUAWLRL1E6UtjAs/MXBOxlp92vha1tRhbI369dz/MDfhB+io4YtVRucPofMGA9
Hq6rnh3ks5uq/Vz4nGbFoVkQrk2WfAq0X68m3HNe8w6R70pMqYYAXrIe/m9lWKff
SRNGmUzPqLsRC4vMoZ3+rYtpx/5lttjGf7CBP/9QRGeo4K8L6rg5agMkuPT8p2zS
aGExPlKGTB2HXP4KQPZ/kwQ0Of5/PFv08PtziuaUpJU6cnq/L6n7P4c67dZLQrxi
lhijbAQ0eDRDI/Xu50x+HUbm3qKkRg8NMsZlnYCSx3a4Jm5fKCy4rCUmHb4/Wurd
wOkDOoJM7G9agRKB++ztG8MwasftH1pT+s/RJ8gsee+hLEAwsgaZmojCwiQwckzb
I5HD2Rwe6CI43gyOvKfuKUzdj4/EzE2sglKZJO8VfybCPvXfslBnuLgDFBKlqFqQ
AYGZuDac7vXSJoh7yWl5l886I6qIHElfRrVEk+xMJ1Bwxz/8OXSzQrEjfeDpV3Je
t7ANcmhGfjRI7GhPO81L7oYK9h25DJqIOLymcYyG8FyB3HFeudpLOpmSpDq2hq8n
JTK0giHIVpDEx0v/GLJgrr/bvpHGS8gXmTngrhfcctsLe4FxPmIvLmm450l5gHdJ
7BlQ4IiM/hmmiYGWotjuHYAqbXtZfAsoaeutULYKwkOreWdcBeNdaVnGOmqQVEJA
mQf0UcyYuRrprUygKQxq/P8rGd5W6+Wc5CTcwrqm1nyF55Ip6tW5IHv31m6U/ar9
7A8H2mnfZ+VBTg2rny6GfwR9lrxatZyh/su6p9MHOACvj6vSgueYbulF4uJiY0AI
SSlF5+oPfQ+UGAkmEuvfwZiSuJLZDCBtTZ2RPRAQBJ7RqrKabIUly12ZGxxozTtE
5LAHKXP/N9r44Pe91535l84zLeu+k3d0W6IJpCxQpbTe3FogqVNKCuh6ocR8zqxm
toXa882sKTzJxhKP0gRmq/Tf52WTY2/i/y7VcGMdLj12eqnl3npbEXKrnTvUw8bj
R3DASK3tyQb+HYd8MBLb2M3glv/Nzeskb1qXm5UHC5vv26vFAgFXxnAdLDxw29B0
i2/ia5yvLq344uXSvFsfUxI7KBho0Bc2TCtJ5mblsHIZkymkodrOXxbWewllhozv
+sZt1HuMgFryzY8XXFALeyjP7FjjAcVFAU+kXchSi430J6Z45L+TPA/g6UsJTy1J
LqgIo/yy7L22rO/xZPZSJv5QRTBidph6tdUavThUWd3n3LEXLdRidEwyEiinFC9l
KmyOoIh/qJBQYc2Ih0FsAQVN8TJnhuiwZqrptFolRbtpcE82uGdE8YOr+wutwB2f
EWD5PW1Gt2D+W7GYU6fYTEt731I0e0OYVHjgQuJoLd3helR0J4shu4Z8J2BotujV
WuSLLY7v1JNsD/vMewCOWhMpHS+3SoDXpZX0Z7wZUjO+nInhnNSh/CCnKVvJbR2I
oYyIj/ZATNJAuky4KhWeTrTJX/hVCWyEic57wOWN5f2Bx8ayuuFYJLGWgl7r1917
3AKNWvfa24PqoZ6mamg0XG2SQ7NSn0Jn4SsCTKyTapdgJ3idZ6HmCACzAW3gMhrX
KjIkXYxHbLByhoZ+xBMQVhJadoDsqX1JOwT1JvJU/f1HIszHu5kOcq4j67Sm/tpg
dW8RpymMe6x1cpFOu0rb/e1tiIxRJ5WbcCc+iLEPDnjSq732HVnNeFe3ahe0UkUg
sqWtE/RqJxq20XAp30TXoQ22cSLH1N9Pgs029kQndKJ+gm5kjSQFsAlEvpx5YHq0
qjZp2fcDHG7wLHEhopCk6EKPjTBfqLuAPRx8Shlu6Sl+mMn0VQDYim9FJnq3BzFJ
F8Rc14rypPcoJqj9FvVm5eI8KkoiEVtsdcJOUWS5j78vS046bW7u7AFQXwrX4Fu4
wn3NSB0WFKb8ekNYyrf3INnnc2vY5YO8BRJryU9Tz4kjVjUDSrbdga7Hbm7DVLjq
IKOnvdIgjT4PBCeSUj13JiGxXdswINSIDX/QYe+1eZWm1TRiQ6/wNmOASPuG8Asn
DVUtwePOVa4WnHaunjFo/qTKSDwMtLaSNm1cGCnMdYnHJvIB9oZ0Dv9R95yFHgih
ej/+t/moq3d/6hZTQ3TmWlRE0SJfh6e95fbyWJ7VZ+dJSbkDQaxLpEE8a+gFXj6c
c/+kVUdBeJplyisgHKUQ+1ycXB4fVvItLHgHs1hIoOB1MyaPioz4fjlieKyUuWLw
bVz/txYLGYzoO+S3ETa65cABZ/s1285Uh5cUrwaZrudNyhqxala5kuGOHyEoi8j+
ub8lzvJbruftkrY/PksybLY/ZI/cI4+jIOYtbug/+ZaofOo03g9S+azo9ej2JwOw
YT576t/ggxje4d53viiEaiCxeiDJIL+zqbl80JqShZCdQXo+sLVTKA65XIKlpia2
XJPcEY+YYfyUo7kzo0m6KValfDErIVkNj3+qzAmg//gujFohzxbVnZrJaK1RhrKO
ENl95h/ylGyJviItzXPUo7ouuJfM9yiiwuEUwYpllsrsC0x1hIQwfOet7cZmr46C
jCLQbBgTw1YQ7IPChE3DLea5qucsqMYLpG874pPFs4+RdIYg5yZcsh5j1p3XVnGF
zgMdtMl0HuncMbBnWnXAKrArVRX3F9+mrKkx8of3MxruUnZyxwfXHaQL5v0ZBsR8
ZJgHhn3dDt3a4WLekCJAIFGphsOrU74r6i2K71Zm3dK0wP9GQf/GgjP/eqN0h6/U
HrShAbc/HBqaRJyZaOlVAHF5rx1EGWvvwvkapHtcI4wVtZNn5RN9ZkJOlMSDAlZv
MiTWU8onJuVcO4gKm+19uGZ4hJNDZ86lhWl3AIZ5BWiyec7Z3iClxDLMTQsIxGpt
gJ/qgUVwO4WzFhKRBMBeQvKGnv2WbDc6N+Ns33/0ZunXq02tuEHFEIx6JSUFNb7t
YPHMvYS4lVGQldFcBcdrP7bcWLZBMTaXCaAxuFnjJSCOr0Mgt5xo1pz2pyg8+OkR
vNdeTNSfhCT/Sns3qqvYC02lYqWyqv1OFiufrCR+mOc8esisRzuszeYzfufFjkjp
pxJIHt4yB/QMCE5+4YeaAYL20qx5mCWEZj/AtPQjUh2XM7SIhfgCFk5e8on/j9+E
0Gt1eTBTSBI2ItGuMcDM8+WnEjHhZ9GEuo3vKlnHf/QxJBctVYr2g0aMX7hi5SJR
URcN1939em2/uI1mKRnTVtmVV7GRlCvIeL0dV6DyJBpY8ROnaIgAwlrK0uzNN2Xe
yLHKnWNsDuhH4A2+1BrhSkNBHaHEdcWzdvqXCpFIU+Mwf0x81+lo2zJ/J2p4Tovm
D9NbEd+DWBrNa2f7oaU7Q+a6d0absZr3jX/fpqjxFTUT3TaMECMbqZ9GpIHFnuLO
WKN0Whn2IL7jfWsnhEkF8uGnIlmAKZOOouyVcO5ERtIDWrNemoCv+iW3yViIcT4P
izyxWi2Be0Nc0tDS7oaPBVbw4riWhwhvnYjxgCEPUJXRGH8c8lzvBwjhnSThn2zA
WO7eMnwpvi2/wwocN69rU5amrgAyk991NvZkWYY0WRE8Mxl0L65Ot6Y/AIoLwCLx
qGSy3+MuVqUTuVrSil49bsR7zbQu1qVys/FZcQFpUcp350NhXJ3fxWcRlJd4MSUv
I1Exg142c1Bk24xgqf0elYikmL5Z6ABPRNBa1NuX/wXq+3lPbFBQF1n5ySyRAH/Z
UOtQ2AtWQivmhJU7bnDDTJucljVjfn8yp28o8nX7Fe0ibtAxewyKjbTM8ErvfNQh
pR7x2B8Zdxddh5r9DGTZwxIoAxmCTNCOFohOElzp1FRc3MpG0TVue0+z+oPaL5ou
KBH0D8FJVNOSfWNq8yQSWtDiJkcYR4MjnIq0hvnacNISd6BxIfT8rPkVT23MYdQD
Y2tcNAU6gGXU9JfFdHIwMtZ5aonztlwxKzTO2Q/VynfE6Zk4DPNXoC6NPQQDXQ+2
FMNn660LoCyO4upDYOqov1HFiOPuKp3YrnOPzBE+82lUZjY0GbQJsIPAoY8o3bmi
kBq8Mr4kMNmv1EazJR8y9Zp6PwpgiyiBa8rl36kwU6WvozecH75divTrqIWH7qiL
gp781NRqaWMBLgd/0UfW+zEG/vasV33xc+2OU3zDZEUQcOzeL2wyYTC6p9MmWVl0
QmHbxZkyv2+vJNa14n2/LG/ELhEJ4jFiyVZ4M9ezowxl/3Hvit7IBgY5kaGDyVXG
+YdI8Wru1e2hY8bHN1vGMga2fToafS0Z2+bWjAkL7oSbvsLUHXzbbZAaSYVFdWOq
86duSg2uWLpx5D20XxS036/p9dyLM0p1V5HQ27njwQoTdaAHY7UB829r87dDs7B4
VqjS2liwh1FkBW/9PCo25SzkK9g862dWvSS4wdLDa/aQBnWCC7wL93eBlDhFCgX1
AFk1CVTHcZE1vF2SmhmWf0sYGKHYBtuCzC/Q9xG71Wp9IZ/Ei7RWnqsW8JBQMzlT
PSR+yVefMYR1ommyJTjiByvyE4QB5WriQPmMql+EBNP4n59TvOz2xNKKG04QkiyJ
HcphyWGdbcpiZj03ph8vMXgH1w0hJt9+XrvEPGJF9Oh//2ZyWP+3OD5kX8Sjh4V8
3rd4E91YmOLAxMVr39CuTz5Q9Dhx9zspN5CKMlqqAmUR11rvGQ88bHO1wboXDKEZ
pMaL33EAxX9T9zaDY7KQdumZr4xc8cnBW6mThSclFhPN9tRJzpKWWk/DC/p2fClB
qdbYRynQf8waxPLiI9GIk8sWpoKjwuU+Bcq2oAJDxseO5u4cOyPWiIBFSHaEP8dg
6DIvMcm7tZAQL1PZhYas8eOmcsT8fxn+qCXmxTB/9ptOqoKgZhC4LhOCkQy8KEWc
McWxb9xt8aLM0rPlVbsyrRgaon8pN5xvVWQKbWT3WSgGsUkhlarEaugl2vXQXW4l
r2AWvCcguxLFWU1OkGErElb+7KaZMacEwoenbpYV+sKL62fVD4ickNVH2IHL+PJY
LXZKZYiTmJ2sGYBSTi6qSs3jkpKgUO9ZbvsPH/BmMKfBuyPcr4tKOZXj9fjEXrBc
fezxSXG9ah58Fxm18thSqQojcmmP/ri+ICdvhBosd3xuU7izbzmbAKZp9CwJA5gj
/Rve/qxKQq9serxwcXhj4YW3wfB8Dqdi/zcehxso1ainWBXiK6EWXW8vLTgggGTG
e+PLL4mi/agAWMwN2XhklC3JUwBCNOHR11BePzDv7rH0Aqf5ojIhcy0CbX0D61EF
fSM5LvgZjDPpSiwZ7MZ5xGW/lox4IEaT0pvDX7gFtd98SId6Qy2ux2jW2yq1VVK3
PFh6BZDBUrgqmxqNLa9mi/4aHWp8EhbYYpgjEGARyIKCrBw+mB0s2eH+fU3z5TBv
+knQynfMg5NfRkJAH9uDws95+Rzg//MLiiInk/yz3JbRSXG4CRZf1DBBwMsN4Wlv
fMZBNKqU5zhVjf9MR3plbLtM7Y/QGj3DG8Zwpe77c2srpDQSLMbRTP6uOcjAtUCL
H7pOx16rVBE9uKKVnuDCu0QUj3QjjbwxPAh+X6FvPQ7tg56lyVAMA17hVdYLS7BV
yKmkl7Ug9kwkMqD50t5z5JKLP0i80s7eviVQpgiInSGVpbqU1f/9sCO1UTdEVBR1
npJWjWS60wE/kBSzJCLibZJ89CP42xqHdPU9Ov0kB4Dvnp511mOw7GOK80sx8zBV
C3loy9MXbWp/S1Uy/oX838yhq/t0kncNrZtyWM/eN1DY9jPWZspvT14cUj+5uQMI
PLDzdIYO1vqhIV7M2ZHEAAFtZ+uf44NKS7xoWiM6zbeAOkioBE6IsuzezGLfpHd8
F+gJ1ow+5j7/8znhnjG9oMulfA9uGMvxm1iUbPVBIBkAj8bwZyeWLrBYLhMBtCnf
Xbvyr5vN2mD8F0MizAS+rkguFJ9f/E7LaEh9RT4Zh8ZfY0QOO1xQXveywdEwSjMl
yfaMfE9VS0Kru77Gw6CA8wa6dt7ZD2e4K/DpNzPoZOqdlc1DLlIQv1T5dtkOAmST
Gz/pIZXz1AGnuWBE+WP5w0brE4ouk0kKfydSw8zE4PeAatSUTejY00z6ynsQITlC
AOjwxE+H2q9HlE/AT6EhnQLbduObAy1U6O8jogVnQEyLcyYdW4ZeYX+svc6ztGJZ
bFkCW/LQ4VsCl3Rnu9HSn4pGUqmcFNL6F/6fJte2T6REX66LEuGP6j7gwe3qE95F
NfLXe+8gFt/oMGPRhZbTcthXuhFBQE2mIYQboUC2cZJoI1iA1t078QVglKKKdBrC
gYSc2c+7M+EEbDogPUGnwaBgtQqbgHT+qiBccSlFURXzcUIPXTzg5LQP3CNz6p68
KbEHHjXiw2RjVfswd0BihGXZbYAZOAXofUKgzJdG6Zq7NvcDyd+F1xvbTMzgV4IA
ZJJ2zYkfGJiJ6MggLF+DjeQbxEwQ3dh49bZEkY7p5YCKhDCCJE1MU1AV0xN4aLPh
L9hJFD6HflSJ+8oWkYc3j4VZL3vsIgVR/NzGzvOJzC/2AMZ4qOCjUkBgLvf1+KXu
XKcJEl6qe4kghDQl4FGosqnGkphoYczalKOm2ptmp7M=
//pragma protect end_data_block
//pragma protect digest_block
FEUHBDdkkAczivQsdg1s1BRPAWs=
//pragma protect end_digest_block
//pragma protect end_protected
